PK   �yDY�#UםN  2�    cirkitFile.json�}ݓ�����{���7��:�{vx7����֝F=�j�wo�����]RWf2Y �u�����A ���w����������?���>�� ���_��������~���������_�r�ï����~U�8�C����ä�sà��Y�Tꇨ\2��lr���^����Oﮧ d
�����!c�R��6S������������������㇧�R����M�8��{G��旇�D��� '}��r�/��?���ç���}�`�T��U.�A%3�����|7f)��d����7d�>�G2�H�������Wl�@������MbG>i�s���S5�]A7,�nY�Id���J"�����8M"`��'���f��ɓ��
P�tяͨ�Z���T7�W�M�OѴ�ؒM�P�P�;@7�f/�&@5w �'�(�<�z�{���qe4��4@e���]4��� @]é��=
��1tk�L"�ptTժ0���"�V8yr�ʝ�is� +�<9��bj&Kׅ���{_����(7�K:&o�D���d15�5��e�&���,�	Pm.K`��2��e�&M�a���w�T�ּ�=����Z�ҭ2���nm�Id��2���~W@&�Q�OO2���~�Id�s�LB�;�aD&�Q���$2
��F&�Q�u'�DFAם�U��)���6j�&�r8ն1����$��j����j��ށ��ƶ��ƕ�vPi4��яz�&u�	�5�D�$Q�@����-����^ż
���Tg�V����&�-}�G�DFA?*�$��N?*�$2
�QA&q�5&Z�4'�'a���T���*�+A�D�3i2q��]�����T皠lhZ��nS�d��^z�KCOwU<��"��(���DFA?�$�}��?d��!��(�����Mo�F����ZP����l����ێ�FQ،�Fb��%��f�4}-6NR$*��d*���_$*��^$*��8\$�jd��'��΍�}�����7�Ɔ���"�_w5�>Ы0BȽSP�����R?�.L�C��CF�G����k��V�QB�6��Muk����=�9���g[=93EՍ.�>^�δJ��x?�ܽʹ�0�)�t�X��b��A7�If�����b2da�:��m�RHQ��Eg�䇾�
KC\�����V�c��L�r���,s��M��
�cyN]g{�fq&UD��3�b:e����������q�1��=/wH*��SI�hR���m�Vw���]6�8�u�6�wvj��G��&��tӃLb;���n}l�BcQ�폭Xh,
��� ,O8y���E�Ր
,��f�,4�
���*�C\�����P��IZ�G�U�ਲ਼�bn��.*�*[u~����B?~�5����\�h!<�]^M��c�,'F��0lG=R��:1XN��'��v�a;ꉐ�v։nb����.���X1[��/O�Ec����~�7���-��1��k�E� ���D!b��������r������w��w����oxy��������w��w���E��%�38�ֹ�rnD�e�QxTCX=<X�=�s����0�f|����8_f��_��g����!Η�;��w�r��G��խ��2%�z��,Dn{F8,��qz@�0O�<W0�=fW�0�+)w�������f|%�3��]>^|���$b��k����e� �w��g�++�S�]����bv���Ƌ��-S+��Ɨa�������~f��0{~���_�_��?��1^|���2q��ŗ3Tg�wz��^DmIuU癴���pX6��:=`�^�\Ƽ��=?^|���$Nc���ǋ��m��c��x�3��6�9��Ս0�L��¿��ϫ2�����-�Gd�ev�x�3�e�>��jp(�緜=�3{~�������JDf�1?���f|%#3���'^|���d�d���Ë�񕜙��c�~x�3��퓙��/>`�W����1{?���_ɰ��?�+^|����e����񕬶��c�?x�3������f1���J:`f�1����_�F��?f��0�+��������f|%33���^|�����f��������׼����/>`�W�v3�������J�qf�1����_�u��?f��0�+i֙�����f|%M;3�6BÎ�$�;7��2�-O,^G�[�̮�rz|�X����xfׇ0�+5 �������f|�z3��]^|����]��_`v}x�3�R1��̮/>`�Wj]0�����;�w�$��ϳS5-i����v�g5>�}�[�`�y�؃���v�"8�}����PŎ(w�|�G�ۊC�J�}��ѡk��P�iC%~��h��C�.=*�7�u�
���M�<*�9mh���6B�T�Fe��]S�T���k��o�64Q9�r0D�`X��/�(SI���r���ܷ��F��5����6R�P�f*ȑ�z��O�Z)�*�HuKấ-�udEr��ё'��2�בM�di�Q�^����d3�����#�ס6qd�<�#k	q�2Q�^���Җ4�7���\�)W���뤡Ÿ�+�&�u�}��5YU��ȒxR��B�c3�!�����T7d�M�OѴ��θ~E�Ԫ���^e<v��nG�^�<v��nÌn��׬��=�3}�K�V�c�:7�K:&��/y�m͐B�N]wS�:���u75�C�N]wS��6��=��S�b�'�c�W>`�m�w#y�kSGN]v�̩�^�n����^���|��AEk w�:]���V�����7^GQ��T���%T���(�{�uս~��^�Fu�_���_GQ�믣8���Q�6^Gq����(7|�]�:hM�mC��P�iP1d"i};پt�����uי��^�=�{����D��w=�{}ף��w=�{}��Ć*vD������D��������'c�Ϯ��W�u��5&�ơ�cc�"�P�7����|L��c�o�ӝ���]�龱�1�7v=��ƮG�U�r���Q������Q�벇�e�ڽ8�l�1��($T��n�P��� Y$��F�a#
	��5W5z����46��($d6��n������6.j��P�����i������������^O�����>��:`�84&B'�ǃ���I� b"T��gB�o���1*��3�����#&B�X�<�v"�vp#Q�B�B(N��!j���&�i�!�\�^�cC\�t"�4��3!��'];Mڤ��"5�n>�ͦ��MqsQ�'�	���7�q�E���t�pQ:��q�݉Rh�	Dl*�L�:O�Ħğ)%t�1%6L/��;�����Mq��!��k��:[�)q�;�g���qæǹ(���>L��(���1�-\�N�Ę�.J�����5�;8Y��k���3�䵶-�?S�����8�%�}��G�I'B)7�L�q�%b�}g���L�c�Y6=�E�{a�Ħ�-�u
�R���R��R<��R���R��R8�۽�c�ǹ(��l����c��ϔ�.F2&6=�L��^pDLlz�����$Lg�t���i�6�c��\�Jbo6Llzܳ�q.J%5&6=����g���r�-�M�{�巜)����<��&�=���U<�=���8��Q���lz��R����`Φ���T2T�aڧ���v���O��a⊐��a⊐��Vm��D"b"�Wā��&����&����&��`���h��D'AaB�L�S1!6��E	W��Ħ��@XLl���Ħ��F�I2�qE,�<&6��Ă���I�����S=�*_�[���%��
V̓�Se�VX����yR}v��|����J�k�D�:�6��W	� �5�5��{3U��"XAk��D�u^a���XAk�1E�:/��	� �5{�"|����V���}��K��p@+�`����c�T�	����ł_:1Hx1����,'o��.	OdЂ�r&�ۥ7���Km�ӓ��ңaa���%���M��v�հ��H���U�,���DЂ�rW,#�2��Z�A[���ᭌ7&�dЖo�ex+㑉����f�Jx: �dЖo�ed^�D��Z&��eF�/A2h�7�"6����V�r��䭌_fd�2� ���0���˘Z�A[r1��v�鰜e2�c"hKN	}+㗉��%7�����e"hAm��!�[�L-Ƞ-�Jdx+㗉��%�L`��{�Z�A[r���V&JQ-��ea��{����DЂڒ�G��2~�
Zn�����ˬ�_&�dЖ�J2��y/A2hK�(���e"hAm�u%�[�L-Ƞ-9�dx+㗉��%��oe�2� ���P᭓��DЂڒN��2�e"hAm�i'�[�L-Ƞ-��dx+㗉��%Ǡo��$���DЖ\�2����DЂڒ�Q��2~�Z�A[rW��V�/A2hKN���e"hAm�%*�[�L-Ƞ-9QEx�e�2� ���v�ᭌ_&�dЖ�2����DЂڒkW��2~�Z�A[r��V�/A2hK�c���1���5�,L��c�2~�
Zn�����˼�_&�dЖ��2����DЂڒ\��2~�Z�A[r���6��e"hAm��.�[�L-Ƞ-9�ex+㗉�����_>����5��e\��6�4�Q���i�c-��A*�\��T��R�'|�J%�A*����T���RI�~�J%��A*�d�G��Ixy���\�(���F�&�� 7�k�����Z��dxd�\0�5�QȜ���ZOE��� 42/x�.
��"]z�En���7���B��`����b�#ŵ��G�TJC%s��0���Ll���U7�l����ԙVi7���������Tj?����M�ꮷ��fp�u	Tl���坝�>�/���F@Qٝ���[#�f|�k�����Jc���hR��_�hkO����EewF)66Nä�Z�Q��N�~�;h���/e������PT�gԙ4��M׏Ŷ�*�]ntc�d�`���� EeF*�3
���bTu�\��6�U�\t�N~軳�Q?lQTvg���;#=��S�ҹ�������kl�.�E��}��������U!�Tg젦ǐ�Iw���E��a���ȇ0����w1�-x��|�A��ڲG_�hˊFQٝ�����،jH���v��Lʴ��)����>�(TN3J0�#Py9a���*'1�ф~�Jׅ
cM��r/Ҫv��u#��c�y{�5��uEvQT^|@?�D��l<g�`[�<�d�q�J�`�T���q1e�`Ƙ�����n<�K;����қا��CQy��8��J�����w��*3
}�w_T�2w�NE&e��&$06��/��;�]KEe��Ee��Ee��BQ�u�PTv�,��/��/��1	/����x����o�h�Q2��Ak���
�!����c�VG�N�o������:���.���*���.�
��j�]-����ePTv�Nꘄ�Gz������k�}	֓1�gW��ق��U���u���1��;��u�P�_&��U�P�_$�5��2*�ZCe_�`��k��1	/��"����"��̮Oйl���}*׀Sm�j�L*���-��-��i�������.Sl�K��U�Ʃ�TO��m�`��`��vF(*��~�j��(*�3��v4*)�!6�ƣ��؍~���5�۟��iF�w�����4�8�r}�+SR�k���ia��M���E��U��x��������O��x�ï�Ⱦ*~��*�>�_�ۏ��%\��w"&Bϻ�!}�/X1�'[�!}�{X1�'�!}��X1�'ێ!}�Y1��6'�����|j�Mo��梤�MkLl�ؔ7%�l��`b������(��`BLl:ؔ8%��ȃ�M�6=�EI?`�`⳿�p6=n��8%�gʃ�M�6=�EI?G��`b��M�sQ�ϱ�<����a��\�J�6w�M�[6=�E���g��w��w�¦�-��T�ab��M�sQ*y��0��q˦ǹ(���l����c��\�J�a6Llzܱ�q.J%�-&�;q�Kq6=���8����wlz��R�wɆ�M�;6=�E��Wd{�a��M�sQ*���0��qϦǹ(��ql��^7��7���g��\�J�/6Llzܳ�q.J%�&6=��8��ǈ�lzAi�m�ۡQah:�T������s}��;T\�&��h��HDL�0qEHDl��d"1��!1��!1��!1��!1��!1��!1B�aU$���S�lz��Ħ��@XLl���Ħ��@XLl���T�t<��"g)7��ԏTA+�`�k-��E�RH`�ٖ��"U)$������uQ>��XAk�kD��(��	� �5{g"|]��`�V��}L�.JF�p@+�`͞�_�"X8 �D�f_���R,��
"X���N7UF�J`���E�1��DЂ�r�$�[!�K���@���K-Ƞ-wz2���DЂ�r7)�[L-Ƞ-w�2����DЂ�rW,�[OL-Ƞ-����V�A2h�7�2����DЂ��m�oe�2� ��|�-� 㗉���[s���e"hAm�f^��B/bBOb2~���ˌ�_&�dЖ2����DЂڒ�A��2~�Z�A[rJ��V�/A2hKn���e"hAm��!�[�L-Ƞ-�Jdx+㗉��%�L`��_&�dЖ�12����DЂڒG��2~�Z�A[r���V(ZQ(\Q�/�2~����DЂڒ[I��2~�Z�A[rD��V�/A2hK�+���e"hAm��%�[�L-Ƞ-��dx+㗉��%��o��_&�dЖ\p2����DЂڒ�N��2~�Z�A[r���V�/A2hK�A�
}I&�)��_�d�2'㗉��%�oe�2� ��䮔ᭌ_&�dЖ�2����DЂڒKT��2~�Z�A[r������e"hAm��*�[�L-Ƞ-9jex+㗉��%׮oe�2� ����ᭌ_&�dЖ��2���!��C�/�2~����DЂڒ�Z��2~�Z�A[rj��V�/A2hKnp���e"hAm�q.�� 㗉��%W�oe�2� ��䜗ᭌ_&�ph���y�4~z�אb��qaP�۠� F�.6� ���|��Tr�R�N|�J%��A*���Tr��Rɲ{�J%��A*�|��Tr��:&���Zr�dx䷖��(	�%�>J�G�keޏ���Z1��d�t0�ת�%�#ŵZ�G��Hq�b�Q2<R\�K��Ll���U7�l����ԙVi7������]FQ�aӷ��m���r]۫lsyg��=�2BQٝ�����q�1�m�N�KH*��^�:��8mz�����EewF)66Nä�Z�Q��N�~�;h���ղO���EeF�Ic�;�t�Xl{�b��A7�If�G�CeF*�3
���bTu�\��6�U�\t�N~������Ee�p�R�)S��XVzP	|Y��56D���0T��k����� �
#��_����R?�. 4����0Tvg�CF�G廘π�ju>� ��Om٣�5BQٝ�����،jH���v��Lʴ��)��[�a���
όvmĮ=ƚ���^�U혹�FpI��������._PTv����˗6��=����bʚ��1�++k�ݸ��]�����Ee�/�o��k���@��ԩ�¤��ڄ��9�T��
�EP��ˮ�����i���:Z(*�~�ʮ�����eᤎIxy�w��G�G~�o�pdv%���tMo�CN9���2�4���l�a���J*�����i����H(*<k��ePTv��ʮ�AQ��28�c^���282<�epd�%XO�@�]Y�g��Vu#4jL֍C��� �PT��	Ce�0T�W	Ce�0Tx�h_�`��k�}-����ePR�$�<ҋ�2(2<��2(2�<A�z������\N�m�i:0�<��[V��uBQ�]��B�߫��S٩�Tg�V����&�-�A�Z���;����mG�2�b�o<�I���G=]���(*�3BQ�I���0(�7�r0%չ&(���۔~:�����]���̓x���x�a�ϻL|w������_>��8��t��8��w?��#�1�� �ӻ뇆��m�`
�Wƻ����1��f
�iG���;O��6F���M��'���V�F�f�HC���q��,)j�24NN��H��N�?Rm�L�]U-��ft���|�]7��4alh�c��)�c��^��P�縇Y���=��e�]S^e�&��������5q��j���|K���A���8���(g����JM�r�U]�+!0�*f����U��� ]]k�R!]]kd0a�*:T�52��`�V�82ڊ0t�EIX�Ȩ9��Ms<ICWq7�~̀%%]��ȘO���ͅR�$	��C&�ÑAp"6)2�O���o�^�=���=����ªVA~�G|��k��ݵ��2M�wIl�YoU�vC�������w�ѽ��{�|����D��AEc��FCS��p����<
>�z���S���G�>���M���D��v��Rl�t}�������|*���c��l
j���'�<��\�����L�?����Ш04�]��~P`�p}���;U�)����V�y9(38�VTfp�u0��ǻ׷<���OF��WG^
����y-L��n��Mw1-38��!~:��W�w�+���i<��O���$�;�\ht�U9��W����x
�+��+�#�{��{�೩�Y��z:�,��$��*�p��W���e���T8��3?'12'�����`��՛Z��41�>|!?8��^}�C~�L���� ��#�o���i���Zq��F�q����;;��ѫ�G~O��w�g���Z���E��#g�؜��'0���������}o<k
1�ǥ+t|:�6�s�����`| JΖ�v���=^��>�]Q	j�7W��'��g]*Q�
8�;���gMwe�Axg�$;sϜ������[:�{�k�
H��6$盙3h��mՔ��\�x�$e��a0��{�ýF]+�� �KE�(.�
�r�
�<ǈf�qNf�0w�u+��3�
8|�0�~��l��id������5�	��#�[rG���9v	-Y��#8ʀ�#.vx��g��[ �Z��L%�hR�I:�<��KmlS�(ך�0�Xת��Ў~��ed<�"��\C`�����N�z55M��;����W�)��L>n]3�����+߆�f���{ƨ���mU4�Uc�N��!5vAz:��u�����7���2M#��
�,3�ܠb�m������C��QH��D�id�..6l,2)������v��R\4�Y^�����6�F�(T�4����SdB1ҥN�I�h��Y~:�-{~��q�o?k9�~�8����lx�TF'! �3�C �5;AXM���E�*���m�P2�ԙ����y��yp�Lo�n����������hb����Q���-q=�������H2�!C��o�m�])�%��=)‸Q~F�4jK@��@N����)c�&��$�܄p����n�Fr�m�In��7I*��)o�[r�7I1I�,~I-���7�;��~L�;n�������(�J�������i��*���r�l���{��H�IG@͘Iߍ�ę��(z�q�4�����M�m/�v��o�[�n#QSl��j�G�eBŋFbg�V���!M}�۽���`�=�n����@�m�IT��Z���p���+n��5C�\5����ذ��n�2VR$��c%1`�J�6��$��d%���*+�9�L�PT&*)���zS�����VԂ�6��Z m��������������/i�s${�+��P���t�kw�O���e@Pa6G-��56O����΃ZJxd��M�y�Bp�'i�*�P��7�R,7�k�=7��a�%w3�B�yX)=����t�C��D��0�V�Y7�>�1T�a@A/سmIߦn�$l�I�*>���m��X�G��Ā6b1`k�l��7���ߦ�?��۞�
D��f%�� ���� !V']l�"QN��$A����A\W�����(���('����֞��a����2WZ���X�X���*��K,��!��b���#����7�í�2�A0g��`��D�P�i���Q�&:��Mt��� �8m��Q5':zQ':zm':z���ǖ�1r7����e�$��a��.��֞�Ju,F	�b	c��ł��d&��Y<R�]@��W�u�x$���5.�䢒�����v�ݸ���]���I��<;�P�T����AeH��7VL���x�i�YP]}��=2�"���v���ȃ�� ���]�a��}9�����(��r�<+�]��u�rJl����"�[<(���ZX�t�ߢ�"s�E��檋<�@��y�k0��.����]��waF�;!���<Ae�� ;��2�(�] ��G��H��WR�a��&-���%âT���N�o�2T�乖e(�I_LK�P����/ɹ䮑���T���f�U��-*���o@�ǻ�~0r�����^bzpb�
�����L�c #�+UPo_5�ʔ�{w>A��#%�oPW�}y��{[�ʧ8H����ߚ%[���Ɯ���|��|���t@�*��Uz�pԲ���/)p�
曀ޢ��&���gN_2����eb�nN_�"� ޢ�9G���.���������i������y�����/��~�\��L��z<I�MEFA&Qr>�Q�I�����?����
E�]k�s^P$����Z,�M=}5�T5+�$��
KP��3HPT� DP�*.A_(ӂ�#MV(j"�@/A�^�a��&r8T>���O��K�":2��wQEL��wI�_aa��-q#��t��mKu_�ڃ�Š�aE�Ã�A�Ê�'O�r:���b�Y��Dl����|q�E+$5qCß�0g ��.�-�8�4N�.�<5�Ɋ���ĥ��$��5������7+J�xD�oV�>Ѿ0J߬��D��2���-Otj튖'����O�a?�VHj�>�g �F��p�id�8t�-O��q0�q:���Aq�id��NC�;�L��q0ܫ�id65�F���O�4ty���X�H�^�3�W���=��5��u+F4�j�1(_�4�=шv��NC���8t�g��t�.��8}��}W�T�_�KR�Ϡ����%�	+$=�O�ϛv�_���r��L���N#�`P�t�j�����A5�i�*��q0���`&o�@��b)����v��vÊl�dHdρ>Ddۡ<Hd۱;Hd��:��L�[˚��uB��_q��:����A����؉���`P���3X�v3v��A����e
�^��!�bP�+�1dXM�^��^�R_�3���]|TE�>0���i�ى�ٹ�K��af��f�#�:�����cq1C�j��kw���2��.2�mx@ΐ���<�V[�N��āD�E3xf�����������̿��?^|��/����k��ǋ��e7��������E�a������KR�	v.�R��c1�?�^GcYW�� K�}!^��7�r���ÅKA�2��Ì�\�q�p�8P����0#�,!��Å?0s7�E_�/S�o&H/]��� �>��� v�tG̀�,�s�<��a�����~3B�FX>��!��Ì��/]�y��P 7B�FxY���r}��G�JN7�e�::�]�y5/���]f��*U�_P��k�9�����n�p{@��a�М���8���eym.|���D-������Q�?.<�C�ʓ����o�̀Krn����7I����3B�FX�>p��bF�K�
� �Wf�����4wB�4�8��L� ����vy�7�e����'4�<,e�n���,�d�= f��������!��3B�FX��p�۩aF�Kjnr{1��aI+��Cn/�!p#,)��y���0#n�%�3�Ì��TT�<�~�aF�K-nr�-��aI��Cn?�!p#,�˸y�������Z��!�����p�<��S�7Ŏ���~
3B�FXR�q��OaF�K�@nr�)��aIu��C��0#n�%M#7��f��������!����|��<��S�7�����~
3B�FXR�r�p'@K#ʘ�
`*�B�HQܗ�y��ۋaFX2�rK)�Ì����<��b�7Y����^3B�FX�3�0p{1��a�h��Cn/�!p#,٘�y���0#�=���Ͽ<|?=�kH1Fʸ0(�mPi �t�@�e��	E�_$=����`�E�̓�)1�_�<��\�`�E���){��Y ���E{��]x&P�-�B�У��2��QT)]��(��i���h�e�Fz�b��P�-��K��"�Bo)��S�QE�PE~Y��(����G�dF��|l���U7�l~���ԙVi7����W$�"�(r+�C+�E����ou��NA38�*�W����NM��6��~A���En��ie)��q�1�BfYfVH*��p�:��8m�ե�lf9�dQ��M��q&��*׌Z�0t��c�Aӷ��k��h9�dQ�L�3iLy�����`U��"��6���k���Ð;0Y9�dCo���G�)���B�*v.:c'?���dk6�~�(r���!K��2�΍EP���\cCtqHk+K!��,�܁���� �
#������R?�.�)��A�!w`�r������Q�.棫�Z�j��S[���V�	9�dQ��lяͨ�:Sݐi�69?E�vc���5;Cn9Y���r��B��Ő[�P9z�.�PV���/WA�jǼn�tL>����ʮ@�[���D�[�]EPP�VxW�6��=��U�b�
ʌ1�+�)k�ݸ&w�M�"�"w�܊�F!��U%�m��mP��K1u*�0)cm�B	�~������öG�߸2D�߸2D���MQ�7\ST��������'?d�J�֕!� U���ؐ�Z�5�U�O5��>h�T�8�v�};败P�7� �c	P�7V �cP�������Z �C��oh����*�[Z G�*�[Z G`K
�d�١5}6i�nU7B��d�8�zl���!���`�o-���
`�o- �?��[Z �K`�oiL�--��� R%pS�PepS�lH����6jʮ�r8ն1������ЮީV\G��7�(�6(�Х��*j�T�6'�ٶU0��h��{�2;Wq�P䖳�՗������m;��������Lj�F?�a蚴vkj+~:����(��q�d�0��M�LIu�	ʆ��)�6%�2;_�_B�[����ۻ�od>�O����~�ü�����]aQ���\X�[�r5T�$��_�l������tMv��:]I�.�NW���������t+|��?=ϝ^�N�;�W�����n�t#�w�Oy0��%��	�n��y�Yt¼�,;!�#�0���N���e'�=��v9�r)��#�n�#�j�#Ə��<e���s8���8�\� Zt�����@h�o�~�*�˳��4>E{�,�}��x��)�k�&U� 7I�S4F�x�{}$�^-�@���Dc*h��1���%[A�d!E�-Ѹ
d�	)�l����
B�X[�	4�w_R���������C�8܏����Ш04Y�t-�N�A�u]>%�{w*N���=�?%���"_�)��P'JL�Q��B�v�-%H�E`�>ҺS�k��xJ�%P�QI	��D�Qb\)q����W}��/�]��F����l"�N�Lmd 	�Y�o�fm#Cih�V����`�fP��F��� ��$P3���h4@kKV����l4@kKV3���p4@aP��F��� ��XC�C��3$<D	ZY/S;7�Qm$<~��^*��'弮`!����,\$Q �-��^"�D�Ԋ{��Dkj��e��S�p6M
W��D���q���b}�yQ�j�k<��C3�Wn��"�lRX
� ���R�����K��ly�v��!hF��������V����yI��2#1p�N�&">˩h���&�[$4	\ᠣY��8hW�BG;M��Xizf!�4YH�!\�i�.��Xj�����k��^9b����I�i��i�+��8E59Q�׵[PdL'��ܳ�l�F�H��w����2^�fV�#-+�Vɭ����T@+���]n#�si�V.�|�r�J�'ؕ'_�/�E��n���`���?��?����<{��)���~s�m���ο��o��L巓ڟ���`��9�f����ov��;�斿��o~�[8�����S��),g��[2L����ǂ�`�u��hp�,�g~��_p�,�g~��_p�,�u�7v��Y����Y���1�d�=��.�n�s�˹����r��<w���=��.�n�s�˹����r~��L/�
s����>�\b�g�+�|��Dh�+`WV�,�v)��,�n)��rn�r���d�;��-y��d�wf�[rŝ��lqg���<��,�n�s�+s?��-���4ݒ�?��K���O��?��/����|�f�����Ձ����p����r�N�`�����_���X��z8���K���Ƕ<#y�\��lV�����yE
���\����.��ɴ~�~�<���}z�O�W��x�ե6�ɂr�)�S6���U}���߿�&O2��*���|��O�������S�����_��������X>��"�=�O>�����q��*�S	�ǔw�Wfd���������toU6|�rC���6^Y�i�]ڝΆ�@�m|�|	��}������?B}������C��>��;q����_&�cc����nx�z��*�������f�^����z;����Ui���t�̭�q�n�Y��K������_U0��k��J;Ӽ�W��Ι�}T�>�o^�[���E�W ^�sPY[}I��@���	�luԵvk�Xk�ƕ�v���$�5)Xi�����_��fYDb�Y�#�YVw����z��/X�*��L���Z��浖������^�j��O'��?<��ӗ���W�w���r@�de���[��˞KYt��|�>k��Z)'�{BP�ɭ�dT�D���y7F���G)e�'�s��q��j9Ki��5oR�W)6������\���L�.KG|a�,��Q�t�|q�<�0��p�dрq�����9��t���)�Zԇ�X[���!�?����d�݄a��~1l�a���_3q=�\��B�4l)�z/X[��k1�Fb�K���}>�_���^j38�Iơ>?�8�^s&��&Nl7/#�0ԧ���^�����s��_�6�q�������~^I��Fe@��0�m����ݏ`������A�%+Ӭy��j�f�Y�3�<�3g<+����������Kv?��\�ϻ��T�S8�[~~z��p|j..��������'{z�����S�C���y��>��L����?���������������������e�+�s�����O_�ǭ�_7���C;=~�������>�gT����O����L֮�}�!c̊�3c�'PM���}�m���iS���n3bl���ÿ�e��R8m5�˾;�!KUp��x��Wj�4ɔ=�l>7�� ������g�;N����+�+g@�g�����E���)w/rZq�^~�:����o��oƝE�� |���/��wu'��wu�颻TwAD�P�}��3���E�5˟�Y��O�R�%y���K1��_��������o�����?���������ӟ~�O��>~a���d�<+���y��y�$g�y��(F�Mf7�ʷ�8������k ��!�E!L�`Ob��Gx������<���j���{��z�^�����7�x�)���Q�o���S�l��S�>�f�W�D�hxݫ�/���l�6[h��
Եf+�]k�®�f+_i��dk���w]q]�:B�9�EW�h	T�7��xv��h�I�ܫ����O'1}�7ν����3�yk�%p/��J�y_.���w��������o�2�J��k��Lo��kά����k��,�Z�+/0���������yo�,����Ԋ�-���A�|�e�]����IH�Z/x��m_mi�.�H|�S|�]�«�������/�x\��fk#��[C��ne�+�Vy��n��k�Vn��b��w�N����/D�)"�oA_�z:5D?d�h�+�A�n�F��Ә�^�6��*�'bK���=є��ǲ�_��Ο�_~��,���x��z���J���ş��?����{P�]1�U�Wy�U�?���">Yt�>o�`��D��.�B6;�4�dP�c��-D�j=��\�􈋞�d�E�)��8N���O����U~i�{B�n�W%T��˧�d�<=���.�����-����ў����ax�K��]:��e<�������y�����5!/L������������������m��%l��?g|x�����oM�h�|���٢i�������OW��t'j�a�*M���c��aŖ	��_>|z�c����_���?ߕ�?L,?���N�\���˿/C�g���ŻS�pU��^?�~m��fM�7��o��[��K)*��ޱJQDI.�3�E��wP�.��gq�_�_<3���U�H�B:p�.im5[[k�.k]�4M���p���[�Zc��Qeͭ���a���G���ǛU��꫚]���ew�n]v����pʮ�(�ťzg�]���{ UvN"�Y�1�l���-�դm�B`�6@I.�?��V���J��Wu1�6[?I���Fܹ�l�.mٕ��'aJ�p����`�� <��]|�S�"\+��|~��p�.?G��ڲݺ�5�^Y�(Y����5������v�WU���*��lV1��lW�7��&�*k�\�nYCߐ�G�����R�kլ[bss�� UNʢo�&e�jqW>�۫Ek����p�_�~�`��f�|�j�ua��5��U3F&!��۾ջ��цX^SiO4��T��t*�=���6$��/��J�Lh�W|�jqQ��,���Q���VJ�=�fyg��u��u͐�o*,�ba��m8����X��X�,�4���[�������`=(s�f]��[1�����Z�ע�����vx�M�"�z�Vo����e��v����X.��vd}y筐/�vߟ�
m��ڰ<��hX��������}]�J��B���?���Q+��q +��X+7{C��7�hwKa	8WUYPZ��U�u`�����m.�1m���mfW��6ߟ���Z�
�)�zZ�y+�S���[����
Wy\T��AEx�D��r��yTZ	%�
�o��W�at��>J�A*u1�Q_w/����y3d��͗��e7H�5��U�$0�Ư,�YS	���5[���<���������\T�Ї��GE��4ˬYS���{ �����k��+�U��X��@=*V�ϐ*b�SU�?l��=�ũ�nv��_���W:NM�*�8;J�z�WF�,4�z�袙����4AM���yl���K��,\�Ywʋvߝ���K��O(xΥ�X��̚9���e��NZP�������p��x��1k��ºыn8�x��b���u�/x���_*"�}���x~;��k�~#����.[-�D����!��^��J�g��hV�S��od�J�B��ܡ�l��	)�JTH�&��T�"��f����"���W,��'��vߝ���D��u�J�:+B:k���Czl"u�m�.PG���{�/ʡ�I��F�T��~�j��l6��7��FFL����'��+�[\�L���oW&ާ8��h���h�$`�73�j��\B�O��g�0ˁ�L(�^s0�a2��U'�|��z��+)T�J�Q���Ǜ]�"�
߲Y%GH�d[n��ݗ����%4Lf�*ti!|�ϿI_�̮��*l�׵n�·hV;�mFn��=9��

�n��UX�·�J矵����R�l���Ҧ�-�Վ]��"W��Q5M���#W�x�D���a
{�*G��w���&hW���� V���%�̭ZBsqY4��f�<�� ��0K h	���� V���_.� ��[��MqY4[��FznqA~��YA��зKx�Tq���s9�6����\\�jڥ�M]�Y��Y(il8�@%
K%�6�bq�͢AY.�f��қا��ǅw�V@�p9p�J�uwg~уlן��
�e-���T����;�P�)h8�@�����l�kd�X��2�l�Pղٺ�����K�ZOA��3��=լ'�_� �E�S�n��Ζ�8B�o�fK��?��cO��
�i���x�O?��\���c��E`3k�q.�����E`<Q����\��n([9�3��H ,���@'.�#���c?����N��.�߲}���	߸���g9�ix��D`}���67\|û��V�o<��d!2{�n(���� �+Щ�=�}���f7\���uW�P�F��)�<� �d��f73 ��nU��������7<���R̾9��Y��$���CQ�&%�2u�����U�능�7Q=��ܭ������f��#�p��iX��fa�+B}#Ef���/<���n*�U�ֿ��l3d�V�Y��517�PF�d\O�P~�QzެR�t�E�-���
�
4�@��'
T�|3o�nj-�rd3d�S�#o+�����x��ͳ@'
S�����C6����% �[<\D�q���n��8�2�
�*s��l�#�����{Qg'��:5�a݄�p�{���í^�Q��<Q*/�s���X��w�p�;c�V@�S�w�X�3�ozg�:�
:�.�C��+!kp]�����1����4��ߎ"��v<�ط�i�&܏�[�WD#���n��QD�.�?�k��__̛-��n��W�W����k�-(!��\YSo��E�
t�l�����{'���3��q_�a�<$����fH��Z�ߌ�b��>L8=؋�uoy�z�i��t��4yެ\z����T�Zp���V|��ןJ�p�=2KL���u��|_�����:�� �þ�������<̛Uj������) �̏l���3p�mcPMӁI%�b{�~\�NǢ,�����D���f��oޮ���ihٌA,��ƶ�����A��Lj�F?�a��1�ű(«�r>fӳ��K�V�bޮ�e�B,�N�!��-t�񽊙�% cR�m[�o�����ba��P9�f�7�	�-�햅����u1�?$o=%T�����UX����L��Uh�͖b�.�w�nA�}�R풂p�+�X����VpͰ���i��C;\�2��I``�
B%��,^�+�,�&��`�7�r0%չ&(���۔<�� W[�r�$�-�4�/4�1�k2LS��#�|y�[s�v�
�;|=�X������A�V��ބ��lW�����Y\~zw�}����?�O������}>�����n?}i?���Ͽ�\&�S��_���?�������Ӈ�O�����PK   [x�X ���s� �� /   images/14933c3b-4ba2-45e6-999d-97e61a94bbca.png��csfMۅ�ؚL�m��Ęضm'WlOl۶��m�zs?������zwUW��{�u�3\^N   HJ�(  �  h64����|Y�� c'��  ���$Q#�  __�"��n��0��j�d�9��ʁ�F��V�#u7�5�ƣn��50��n�?�cm$�?���.��=~����t��&a�̀����3x��e#d���I��H��+j��ʼ�W���\������U�|Y����1J���0j<K��=���&�9�7����<��K�QA��-B!�[d��p�+e�c�n����뀿��T��!?d�� *8�[����_q?��LPW��'���Yx�w`W��X��ꈴw~��E��m6�Q��V�ņ�Wߌ�m����x(≥��\�Q3����ʻ�ӌ��f�p	v�AU�rn���ŷ�%�1�)���'��%a�sO��U���rӶӹ�p��"��w�ʽױ�{xj�㋼4�(��4���n��c�7eu�P�K��p���hv��{�Z�����q'���20}�_gk�3�F'9_����.*[G�6��j)IH9�X|nR�:�?��0!�@��G���B��i��M�R '	3���Elh�X]	�qӢ�����+����&jqy(>��=���������Ų�1"�����1�~��%�]0���N5>,�Oǩ�K�\���`n �2���P����b��m��[8��X�3��f&8����4]���UH<��xa+������0Ӈ�5e�e�B��Is��>�����AT���W�mK\��}=C��ie�)�>��ee+aM|�i�K=`���OrƵ���O>*$:9ݭ8����)!l��g�S`�:U��j�,�균����o/<KNj܊�}����t��� x[�nɤ�Zr�[a�}{�b�q'(��W���O0z�n�0��� ����tᗵ�B��
4ɑx\�^9"��:}�_��IH:)��۽B�{o:sN��u��XZ:o<��4����׾��I�0�M0���B|�k�y���0��p�<����X?|�g��T����&��9k��}�lb�F����d�t��2�;T��v��C���`U�:�8w[-#O%>��N![��}5O)�e۪�-'f��4*=���ƺ�~O<���X�����(�1T 4p͏���2v�*�icd�x�S�����U���|��k��z���K,�Z�4����q���_�Jqk�������6=��c��{�
=\D�fƃ��p;�u���e<D�$���7��\E� U�6�ll��-l{Y���DG���ц���@�Q�%�o��z�hNOd OlVw\��W*��B��NF�A�~��qv��h�����ĺ�px��L}n^r�>��RC.�֏���l>|�!lZsI?J�rn2||s�jlo:?j|� ��g��2%_��v�|li$(�7�J�\�6���6��z��~�|��n�9��W{_X�J��9����;k����,�Y꼚i�;�؈����s�&5�O��=��L)2dx��ϑv�Kk��+�>!��d��W��?r+����
��L`gQa:a�� SYֵ����b&m�D�0L���V'\D� 7�T|T
����J/����%�'v�xڅQ�G�I��d�"]����}4��}�c�}��X�Ք��(��]�E^�D]��f�V�|a�충g�#��^��F��m�mg��1����Y�G�����}���ږ������˴�'�c7��c�9Ρ��H�����^ T�q�����
�h}�݄ł�j�ȅ�TiT`M�U��&Z��r�;e�1�*��{�^@j�#% �ψ'�$wcT�l�)9,߻��L�'�"i�K�D �Om��ǝ�j�l���r��`��[ru˰|���g����\�Q�y��cQ*
�3�_��V}u�Y������-"��4���������J�h4bb�r������f�-S��e��&�46hW<��u_g�����M!�E5�c)�T�t����NOx.��1�YL��������܂�� ��V(0�6F�
�K�n�Ov/�X�cPCP�rrb�u���[��l����1H;nE?#a��s��*��������q��ULQ-s'������y����rСsr>�B#�uUK��i�}~ֈ�?N�B��πgN�u?dd-"�%���̥��[A6%W	C�	�����Cm�	�/��Ⓨ�Z���5v��#��9�v�7_��&0�i�2b�bNP1��M<`�v%��>�!4~��9|�'�n�p?���T�$k�~�/�Q�L��v���G�� �VK�����e��*�c�S&ډf�Q�F���.��iZ	[������+#���Fn7���|����.��w�^7��ziM@-G�W=�'���D�?�& ,�uMu	�q�v��>}L�|���6\�>z�|��=�Z��݊�����n�?w������m���3�Uv��)3\	���t�՞��Ѥ���d��N$!#��TvO�9�JP����F��E�G��w��V >�!7����y&п똌Ҝ� 1u�v���EDm]qL2Z����揾���3|V�U�m�Ax�ɡZ�<�%�<�R��d۾�b�p���W����*[�4u�S@����Ll;!"H;/��.d���b m���ֽ-*؋��W|9<�cL���A����H�p�v��Qkc��[�t�����4a�n�_.�6k4Ń�6NZ�����w�Ӏ�j�I*��]YD�G ܓȗ�	LO3Z13i�oJA��-�����MX~?7b�aW�u��i:���.��<ls���U����y4���'���B�vy�n��������7�P�bP�3W�}�[�K�-
3G��z�Q���V=��|56-Ż5:�I%D����1�I��Oc;���4����!Մ��a��XBWW��(ˠ�I|�siq��gkcc\KK�R5avV�T����i1B�T�PЎ�Bs���z��ζ����Tp� ��J�|�PK��J�gX1��h'V͞A+	t�u���W�k�ழ~����I�,��%K5��ړ�F�+���U�+���\{٧Y��p�O�����	�F{5⎊sv�gG���э�&�~7���|5zle�k�g$M(�{J��YRu�	F0�d��`5�*n-�.��:]�dY�K�X�`�U�?�B�E�����<��yV�h�U���X���XM�e��dI��rz�����O<$�rjk!���Wi0�1@cu�]*+t�u�x�d8?���؁�Mõ�z�U��w��{1�t�]�؀vC�o���kʒޖY��ԓKOSk��[떸�ʴ�M��$�PH�B��SI��/�<?�޲��w�ƀ����6[�_U�]qk8	���P�wq��k�[��½�Sv7z�Ǟҍ��q��Qp��$���g�d����Y��3u��鱦�4�T��gDY�����nL��cy�Ƥi�C�U��]���2r���1TeeM���G�pz�^i�%o����3ꅣ
��@"�|L�W���E�Q'�f�N����81qpp�}�=u�Y�>�����gq��w]u�d�v�z~}~xs�O�0vi�S��vd�/��xv>mjv��|O[7�̪�!��wE1f�Ē����ڱ<�����*
��+�A�sA�յ����R��Q8��d3!���s?�21"FE,���1����H��FbV�+T�~5��(�^Ey���ў�33B�Js��Єܿ5lR����gw�;N�A�$M0<x���
��4-��Q����Kͦ�ߝ+U���&�m���&R� 3�Ӕ�2�-�.�����W��f���$�"Y������"��݁� =�;��I>�}(F ~�!+$$�c���ʴ�j���u��q��j�p(,//�,oM����oʖ����ߌK��lq�!��"U8��E�C�n�~�B�i,5�z�C��X��m�^��럣`LP���_�%�/��9|ԡ:�v�U�?8qp��BkW���\��e�����>n[Z��5'��S����Ҥ[����.���rqݴ��S��m�?�N�Z-V��:��5`ٓ/�,oA��4���wƨVW:U4����cFk�"ۏ�C1n��y��e�h��Y����t���hs��OEL�����ZRjA)��cӰ�����~�uf$}�[8�T�m��P��>9?g���I {؅F��dm�a�c�4�N[���+�%�|dB��L� �͑u�9f�֝�����Vtr��ӓϣ��4ԁ���o����i)�U��3��*�Z�z�3����U�dǴ	9>4d9֑?�o�L%�ڎ(Z���ɺ����W,�\��Έ�_L��g��/��4�&_�7��ӌ�܀�β�@�a7#+������5�9���7\]]�{���:��|�u���|?_�����^��d֢m�kvޖ�]7���{�|j��<Jx���Q�q�^&���XV�RљH'�)IOCԣm�GdQwE����4�Х`���l�5���s?��2�q��$��w~���5��Xż)~��m�!u8��/$�TFu�qx�o �3�U*D1�jPf�#��Q�"K�<u�߀�q�� �>̮�;�c�u���B�.�4-S�萍
'���ς�c�qvj�vm�aw=��Udnԓ�̈́3)c�D��ڛ�xa�Yq�ŷ��,��n�>u��2ʸ5;IL4�L4�j�9�(-�x^X�l�w�LFDMO���e��&d�6���,�����}J�G�>t�:0jy<���iW��^��pMN�}D�5��S��6r��s�;:�����3i���k#CˉM=��2j�����	��Efv�j�<鸍�O����wX�V/�z��X� �� ʹ��Ҟ�S;�l�.CG^~�m!J�O�V�^��!z���&���H �u�Oz��Z��o�����0�^$�#)�:A�;$����Y��0���8�r��<)���iM�r�S���Ӥ��2}��.x��������
��K�e?���'��Ξ}83^��xz�mga�vj?�F �i�m���o\li+�}�a��^?q�c�uы��>��c| زj��=a<c��T�[���e#1�O���V�X�75gP��b���� �8=;�T	C����f`��;E�S��.�����r.�2N_�6�_�C�_�
�`!}������xR��H�ӂL��gT�b��>.�h���{b�Z��&R1�t�|lso� �?��>��C7*Z�O�p�	.G����a���#L�F��Go˚�:�Y(s�kxXvx]���]����ܦ�!Y~|���{�Xk�YF<�V-�J�*ǉ%&6�i��������mN�'ot�?��5�т��Ƈ��,�^�^�����ٔcImQ�Ah���Qm��0'������Lo!����E����/E}��v�z52%��RS~���g���"G/�j<*<�L#.��䤓���䝴{mja��o�O�n�l5�,ЛB˰�@\i0O��I������h�c x��)��$��\����?���I�vqro�C8�Ä�c�Nf�\��TS�|e�UC��.7�|+|�5
���3E�5�H�I%�"9�N2�j6�zX�lZ}�<�j2m�S�F�����6��'����uT���I�ک�ge��(��1lC��M#C��JN���e�f�_�OJ&���{�韔�Ih���Vc�y��i�ꔀ����I��J=���n�]���ݮ��g�6�Qna}��k��<&����s�د�h�@�Ql���ʼj�9ʍ;I����z;�K�r��F'���;V��,�#�����2��ˎ� �CiA�6D)؟f��FZ���	��'�V����q��\\a�E�9�&T8�_j&�B�����6�^����Q%s�-����e�F�ލH�G���O}�9U3��c���-��չ��`2�<d^�F �L�j���*U>��Y9��� ;�l�8~p�-�^o����F>~3���|8%ι��WW��ҫX�t���%� M��!���J�AZ�(�����0�_sCݩ#��T.QȦ f?�OcUA���Hw+�ι�W����*M��Ad�K���jH~+�aQ�G9f���!��N����D�`���e�Y��|��%�Q�d��
n�>\Y
�J�AY|���]�п�U�_��G����m���kX,���!�{�����&_��@�$�Μ0l�њ��eSS�c�GN���.��!e�~���c�����:��{Q�"��G���V����w�M[���uk:������!�NV>O!k��O�4B)�?���߲?����%�@Jg�����fU�62��(QT�\;�r%���MЉ�P�28[(���-P��S�;����Ȩ��L}i�Y^S�	Ɔ�J$[I�V����+1`�^|� ���L�Lؤ󹬓ެ�	W�?c��g�Oy��Zm¶Nߪ;��wB�BР�����/�Q?΃�J14�5h�~sA���X�
��e��Ƭ{�VT���9����\ƫ#�v�r����_�h�a�7���i�J�ƎE���FU�-�L)�9�
k/�Ǫ�.>�U{�y�� �ޞ� �o>$�����d����P��5K�1g��2ef ��NjE=�
.�5�MIi��ۃ������)��{�CM$;d�}r�@�w���xi�ʂY3�A����@*�#E�"W�&�b5�y��D�f|R�>m��I*{�b\<�]U�*%�VR��bV�g��_x�]k�"�@���@5�� U�q6!+�%	ۧ/,=�D�|�%���z\!_'^4Q�j�>�c%\(����.=�ǡ10�n[ˁss�Oo+�X��f�$hƤ�������U��5��|��M�V7ý�	�p#R?�ߕ���t'!i���p
���u�?G��S���j��S�B�q�zd@�����f[��a�HQb���_C3��'2�����+X���ze�����'$XiK���ďf�a��z-��}&]��ύ��P���~Wb��̓�hT�q�J7#�?'ޒ�'U�x�4lپ�$ʁZ0���<{1Z�z�s~p/o�z���NL!��6��q�\����E�����2 �n|3\d��d��O&��]|�A��Iqο�b��^�u<���"��?f+�h�c0�=Z��]B������9��ٱɎͶ�h�\k�*��?��Kg]~<��w��-�p��~�郘�C���.mêyq'��� �矒~-��<7��#q0���I���*]�a2�����$����T�M��Ha�H}��Ր�WjvL���p15�Ux
���&M~G�칇��Q�(]Q��I(�˴�_y}�[.7�]�D��|�,'�� ��+�}? ���S��=��n��|�L������s4��)�**�����7����ͤvv�����8��f�.��gF�%Nh�,<뤠�%H�J�rH�$d�
�V}��M�+gn����ϣe�ӇW�C�� ��[c���	x'��)�˨\i�հ�=���!M$I.iI���qu��͢����:?B�ͫ�����nt� �ԟ<)��֓�	��(~��.ڿ�^���|ޒL�tmJ��xz�� ^E�� ����zez3!�Sgu�¦4J��Uc��y������cvF��/�_�o|O�kF����)���;��m+9R�I^�Y�Ύ�����~��Q勧�6m'EH����0ޗ���%ن gJ?����<��|���oN2�׭1���cSΥ>fAU�Ϝ��->K�Җ�l��s�~����4�zc�]����o����5������6�Nwqc��a����6�f.P o�E���v�K����{�f�`���*�ϣ7e����Dg��t�]Z�x����ChY�gc�ᶝg��	P+H��p�d�0_��f�ع�k-�H�oŗ_�_�:ʨ���]]��c
Ά���̭d�K�̂(����W�I�d	��*-���W�M¸�޳{�ۊ�3M4j�y
����y�.���\��l��k�i�W�����A��q�BAh芓���.�fq࠰�5�^���0>�F=��5��W���{���ش"s�$*�τ�"�����T�����d8��!������:kW���}��y����ޟ�2�� ,�Ap�[iu4��G`�h�pɨӮ1(!��ф���(�e[��Jx:�H9��Z�U�on����Q��u#O�Y5}���Y�������O|���\xi�2�V�/m�sFg��J��0�8�x(ݾ˶�O��Z�2�oD⽟y��~\Q�}[]�<ݸ�y�8��$���NH?$l���P|�7��U19p���=��)�R��O.��Æ���)��:U���:̨N�g���s��w��!P�o[&Z�Y	V6� �uT6�ϖ�/�p�h"�D�b�q�6t|0ZoG�)H���@�6M�x5eUM�q~X�IrC�J&^���D'w<#q�KZ���1_�ԚMV��{C�3hH��Zޞ�t�>�l�&�x]7ݏL+@@-ɸәt���o���>����O8��PI�B�'	�l~�[ƛ�;6��L�1�,�'y�A�?w)�"���I˟ڑ����f���+Ձރܷ֝}�Ib{u���?��2{��"��7�|�uӡ/B��7������j�z�0����t���9��-�q�}�������i�L��t^^�?���r��zA�7�����&�{����A�RU�nTU%�h����Ϻ�£�Y��̆x{��_R�:!�}\��^�m�ao���ČM��v��<:������i�"�p��	�a��}��`���o�E$�$�T�r=�@�T[Od�ݴ�p/z�����:�1�roMR;Hj8&*���>�/ѹ�`�>��s�X������l����r�@Z�fռ�w9��铮�E=ѥ=�d��}��@U�F���W:5����#���t[���FJ��KKz�/V��}�T�҉PO[��	�A����9B��ղϩ0x�_0Sr����K��!��4Q�jeN���7U4�o��Y��p�a{=��X�AH����"����?�c�4�>�]90Be�͉S �/�-�x����v�eG��wm�f�w�%J4�⟭��Q$��k΍�P�r�CZ���c���L�m3�1�x��9��t��z/�V� �<�/E�3ly�c�F.�?8	b�}P+�B��M��J+R�
�4��6�=(����@�!%e��+ߴ��s��J@���DwIK��Z��0{Ja��[�,��迷��J�'Q��w��g3c�E�1������I+��ϳ%�7�\P��6q�K�ͫo$�R���^Pdi�*kPQ��l>&�c�CB�*�=���c^�J��5��P�\�
E|	����I�L��<��C$ ��!#�qQ+I�&J�C��4;:��,@��[�7"p+?����!�w{�w��<YV����Q[�@��r�	�Co�W�<�*y�ls�M͢�M%Va��
�~}�q��Љ``�7_}?�8h����'�C)�=R���&O�SۊϞ�	?��������2��2~L/ńT�Y�WΌ{�ɸ���eЉ�E\%q�BA���
,�/��3������K�C��*�fv!̛5r�!��D�/�#�QM�2QX��*3�۹���.����;���dP}_ߴ�M���=���@��_���s��}.�u�$MRdH��>A��ndn6���Q�.���)oF9�o8+���K�H2�Mށ/ވ��tL���ť4��W��q~Lf�E��-8i,�0c����
�2�y}� ��$h�d�Wa�����A��7�!9��jW��ڴ �S�g�L�;���05�{�-��X��#��b��+������ ��
�ԂYv@�q>!�3^�@�U�q(K�a��=�e�1r�&yGr��@�5�c6���p�(�
�ll�u�A��8١�[�?�ZA/6�>�5��Ť���f:E/p��RZ�bGe7���0
r���=~C*�-�^�`EH.񼹴T<��#,�"�p�R foR��a7ty�(�*���+Il�¹o�b��S��f�����l���0jا5��\�J�s2t��H�N�(�/�6�h'~�M��x�u�X�j��W���i7\D	h(�+Z5^����Q�rRE��:�p>q+����E\q��0f,��gG��9� &RP����I���p���{�(}�c�H��ˮ�-� P��H���*ж\";�;�[�(wb�S9�F谽"ݷ�A?�hx4��Ҵ���J~,tM�S����$�K
`�F�X�A���B���m��$M&��,�X��sa9!Ǽn�j		QL�ٓ����w��C2��);;;��{&=���2�﵋`�l�F��U�]�pI�!�f.6L�r'��'��Pۃ �%��)z�|"h`j���B5�����h�-�@����6#hF�G��ʄh�5��q�KL΢S2��1�U�Z�.Z��b����X/�2��a�i�M��^��8`��}Uk��Wg��jU#��#�P5k���p�+1�����h�oy5d珕Q��=��*�/��ZOȍ�wr�+�nD_w��-^C���X����r�ٓ�F���a�U���[^�d�0�E���k�n
�p�j�C���Z�Ժ_a�Z�4t��h6�8��6Yl��>7p�S*�p���G���k$3P&DݦT���z��]���Pe8�Z4�xF7�P'�h�`Zͦ�%�|�����T7���:�V�ˁ"%!  ��UHV 9X~���.����MGP$� ���0���B�b�U����8�)3�-��T�^��5j^\�$ݤC��d�T�v�s
I��`?a0�L��:�f�]�*U�j^��̼ ��㞚f�� �#�[��XE����O8Z.�Z��������!p5��+�%3.�Y���gn�����)�q�n��k>�x����/I�
����e�?����+���C-*�������~p~c?Z���
����-|,�Eü����X��7�v�`�t��6]�/��9V��f��܉�l���t�<T+��Ƌ��&Dɂ����ۋb�G�u�
�؎�hNy�:-->�r��9����װ��N�ςZ��	mJ|ޓ��DA~nmy�M�Mre�S[�o�#+���>���W�I�Y�p<������BK�={�cܯ��(��p��v��%0��c�-Ww��C�A�K��X����́�H���X�5ݤ8�<Hѭ��?]{�t���-�p��v�Ł��9��t�V�� �7�(���FlNFC�2�v�QQm�-�f&��ơ��"vJ�=O=�,�9{gx1igJ ���zƠ�)A7H����d��6�R8�����2b�D�
-�?��Q�3�~��&��g;�XΚ8~�a����(�8�Oc�7h��P�p �ˏ�.D`t9mV���V�� ����A�������F˃o6QՃ���	��t��@b�:~�~�CO�_���:Gz����Ď��������郣O���z��c�m��;��z[ ��n�@�B���sܔc���Y���s���JH^�Yy��l��!t���A���jh�j���JQ��vo��ISTR��_7�}�'g\Bu�y��
�fz�!ڪ�2�l1Tg%��wx �'�T�:  �K��'!�^��֌L���H-V�V�_�F�H	(fFtF����8e1D����6��#�&���<�ޥ/��.����X�-���m�l=�e->^n���i�v������f�_ h�����oAr�=�n��|^xK�J	�?XX<�aL�#�5`�(Ƿk��_��Oo�$���6� ��(� �Jź��U�YU�k=��<~�6I!�kvh=���ӥ\eDx$v���]o*/t����ol���.2���@��U�jm�d�!�ϛgվ�mk}���g���<�у ���q�v{�^#���[���3A���u�_|P��U7� (�m&A\J��5��u`+�..�^̕��S�Ӧg�%;*�4܍�:ձ��� Ȕ�8Kђk*ۿ�wD�bF����¼⠀1G/f��Ŵu
�6uU��)�^��+�+τH�5C������� �_l�4"�㸃�6�Q��V�	wqq�i݆�?];��{ +:t�ږJOo�t�ژ֞��>n3�_2^�zF���N@�U+��8��bV�*�A����d=�@�1��;�.̜��f�9Xd�{�*�:��H�Qg�	Az��6��%h@�?�.VB�$���C����1/I�S$�gf�=
Jr�y���ƞZC�n�\}��1ܓ�
��V�*]��m|V��i�.N�nTT��v�W��&@�ƙ��H� �U�P��Ȥ~�褠6O��km�P �Qm��گ����[�� �����l=ʆ�G�ձZe����b�%36��
u��N��{f,ʍxg$Jc+���+u�
Z�2�b�Z����Gǹ���7�)^ ���)�UG�,�_#V̧�5�ȴ
:U�]%DB�v@��`T��n���ǩM�u~�E���ώ!��ǰ���wؾ�@��{�8I����"�Σn�h��G{��8�O#X�,��&J�t��W�����y1�p	�Q�#��ːF?�6�9Ӈ��"�#D����8�Z�Q����]`��n�
/#f}0N����rب�h���R&�fP�$ ��T7��7[7|�:~�dl���)��T��_"�P�sVL|H	K��ٳzX&�0^���M��0�S_�ް櫧�D*��,��1�E���wj��̈́�>�e)<�I�@��B�����L6����wؑ+�љq	�
�2��mQ}/�7$��G�[0��^��~�kW�#�}8�� :�m� =$�߀>-�k�J!_S�#�h,���wh fL���1αx�lXG3������ҹRֹ�>�����u7G�E�e::���o���u���W/�����	��x���ۅыu�(M�TN��3E��q�qϾ��p��6\р���1�}H��*O_Z ��L�5�ڢ�\��ُy}zL��u�1��b�0�I�8;3��D��n��]}��~�7;HΔf���7�*�=U�W�]
����.���錸�d������g~FK��céը2͂�_Ũ��P߸
 (�!����0���>z�|���=��!�XC�k��f0^�ҳ�I�,���`�5�����[��C]�Ab7�L��'x�jYh�����-7�ӛ%r3�9[�!b�N8M�̫�ؒ���r�������i�Mv�.�Sa@z�!�Q*.V"�N���O�Ѩ��} >�gS�H�r>v�����IR�ӎp��q[W�J�R������UYNO�A+� %��eڱ�3@�1���W�Κ�����VJ��(-�����xD���U������ڃ��l��"N�Fb�_MՌ%v�줄fp9=ĺ��;ed9�l��X��}?!�:�p��0�HQ�� v^�K(e���ᇏ�������Ǎ-���x�96������T0�6v��a�&���j��a${�<�4ן��XK��8��+ȴ�܉4� ]�:��ѻ]���}D�z	[iIۂ���sYhUyY�|;fT�@*�Јѣ�օP�]t�M�'��u.(/\�E���A�/���7p�!�����Y�Z#�CM���ue$�b�X�63up=�b�i4��AY�5��|�9�p��6ēsj}6��z��U�,���;F���0Ǹ��C�9�����ioX�휯��E
˳ML�ï_0.�|�/�M�~���@�	��s��Kpd��"B_pk�j�=8" p�:-�$R�@oG@$�ʚ��U�q9��P�  ��~��hlr4do��R����0V��Q�넯��<�85��wl��`����Ɣ��.���7���s��%EG�ȵ�j�G-�><8��ǂ��ˀE��f�}Mx�}�  Yvj���l�t�4�㠸��}P�U�yk���W�G���E� ��y���Hn�׈����BZ���C�`"*���ϝ)iv�D��v(,]Vt�l�)�n�JQDjBwx��_���<�	#H�nWMQ�=w�}$�� ;�,mR����������w�Y<����,��1�*0J�J��H8P�Ը�Bc!�X�#Q�z�@�>}\�%zǟ�'&q&�t:P��q�*�7�ԠS�lV/3��-�%��.P�����C`��t&/4��i�8Q�P�u.e���u�l��q*8S��z�GY��F1�M���$�&�{�����׊~]�!��|��ou�DF�6�eд�����v��R�3{P�:R�����M;��#H���WXKW����x�1Jԉ< ��=���dm��C�2��U-�+����h=:��N��
'�LQ�/	�'-�~� s�ѣ�k��.�N������C-�����4ʞG+!�5گ��1E.�c�:*�"B��#%�4��=jQ��%�A��n�³�c��/������Xm�MPT�CD?Ȁ����A�k��ʑ���.1�"Q#�
�Y��[�.Ɩ�Ո@	�R��2D���R@9�Zy����F2�DA~�,$�6�c3��촟Z�~��
���d��ㄻ�M՛"�?�~�:�w�b"�x(�$�	������K $���7Zϴ�ynP5�.d�����9�E�0O6i<�����GB{s��cqft���:oa�+B&&��>EJ�A��9���p�,p*�0|��?�ƺ��G��04ɝ�nHG��
�ϐ�[<���Ź�I
�U�5D�k��e���!�����#0���f!P��h�U��K�xTo{����_�m���>Y��v��݉��w;U���Aw�Q����@�{@�@��V�[i��=������q�:�Y(FNM +�مq{+7��_��Q�<���-5?Pa��k�hdv����Q��k���|I��6�� ��TƟ���ؠJ����򹊩�@�L�`�������V�G��]"$�	7-lQ�{q?
ZUβm������רu=�PS�%qs5�?BA�մ$f@�Z�Bq☘4)�:)�sK�0ȝx٘�BY����"T�5#��bDe<�f���]�N� _��1�Ed��=�Τme]��ńV7�	�h�z?d_��t�}r}�~�4@�<�i�t�R7u�
�\��]�F��������P�p�a�1y�'	?���W<��ş�qb�H�~Њ+�#��tf����!�+6��8K�����5vG��L��|S���T,�f=��I|L��u��j.��U	&��5ƛĄ���K�][�L��&���p7$o\�Sc��̸��c�o�P��uy��=��4$i��>z�����^��Itv�6�}�ҿ��/ֿ����d��J�Kq�"K���������F��ݪ��$����2�{�q��~�2Q�=~s�o������ r[�ڥ]�q�X�oG���{e�XNn8M��uJ�?�tcyi�v�oO��¹�z���}��ٔ��V���i��0��i����OhE�b2�9����q<wM�d*J��"W�6L������~��AH���V��7d!S��=\]AlO�|ތ��V�-C~������v1tI�g���m�4,�I_*��DЩ��J>�<����v^�x��k;�a�`m��q�~JQ{/��YX�3�����.�d�)�w�y�m�Y�����n{;ץP/[`*�j�e�[dͬ��n߃�P�I�[��J9ل�"4^�Δ�V1a$~�y:�!tل^�+�G}O�����VBઊ1D��6�<��_�rImjα��Z�6�2���s��d����08�� ������Ao3�xv�g�{���R떩��k�H��<���Uc�*�[��G����mF���T���V��HǮ���]���X�Iۧk��,�D,�����2ӫG���x�f' �{���phRF�纎�V�����4ܣ>�����y�e�%~�h�#J�B��w��dd�$0m/����Q�:~d
|I�ꯘ-%��E(r;{�vϼʹUA�����v2�j�%�tdεrVD}�w\�P��m�O̲9��������+l��4O4����).A�O�ʨ2�d�V�����%���)��͔�@�a��W����V���т������O��J���C@���H�GF�ʰ_����X9�����/� ��,�ݲ�28�yڗ���ř�?���������DEsg��N�9M�Y�l&�VD��Cv�K.�Jl��
�Oei���gK���tS웞�I;���a����Qc��M��ҩ���厛&�
�as?�d���	Nd�N�vi�Y�0��A��J
�?\A'��������;26����;���p�tW�f
o�B&��Dɮ���](����J�-7�)�,]&o��*�Vk�o~Ov��+a �o��Q����*I���W�v+��&9xK% l�L@ �c}�E������N�6���L�a?�P���lU�dǵ�52+�΂p��s���s���f�463�,TX�d��;JA�7��:�y��S˪�eJ:�%e�xf~T�s�/�.7��!_L�b��J�1W��P��o}P����NUdd�!]��$T�����ؾ���[Cz�zd�hU��?}K��/�NB��%-���e3��dGcE<�K]բ��Xq�����
�����6_FY戮Vcx���,>eW�PWؿ���/٫�Vה~�7&ܶ��Y�����~}���v=[4љ��Qe�I����x!��%QU$zaO_ᢉN}�;��2��o�����Gb+N�ͬj�����hM*]�$|�T4��l���X5
r����
ul[!�wr��G�e3��9JqI�&/�@Ǎ��U�Pp��7�3���n��O�Oy�;A�2yb�ؙȚ��� 2��P+/
�L��j���6-����g�QR�����9l=��v o&;�.6�I.�����8��%OB5$��̸ה����s��&�D��bK��$S���ׅI�|�$9��gZ��T#�MC�]�TV;�s��L�2��&j���3�*��%+�
��{�9
�$R� e�p��6�m����,V&9I
,����A�Uw�i��3��Ǚ<�,��C��eoۼ����&����7������c[?l���;�Y���5�-�2�d�'H�z�Y8a�j�)�ЧE��4���(Y�/`p��L�/ۿ߰���|�f�̉�o�ެ���h�8n������*+��`��F
���
��k�S��̪.���O<�-�j4��틚�Bݵ�Z����������D��1�݊��ZU�Vz�)���3}ie̵����Gu�,V�g��:�5s`fE�B$4�^�7� ���<W�9

����?�X*�nAd�W4��l(Qb���Slv�\�G&����D�'�a��d>Ɋ	@���q���X"}��$�π��]#]�i�ifK��zC�jQ�j����/�}��:f�(������Ѱ���4��Fi���n�đzb�H�GN]�fu���~6^�=*�dql`m�N!���ѾS鄓��y��!jՆ��Y�tg�Ս���0�y1�H-g�da<�j�ڵK�0�}CdόH�C6
��8��e���l[�[��%�x���k�a%�7�R*�4�(VaO�x	*y�S#��Jʄ����d'��V�{��} ��%��zRcp ��K��fN~�nҏ�4yPRU#)�4��+�X�ȉ��u���� �v��e�H�i@@�ߋR)�h�a�(���,�T�� h��2��?L"g����y�)8�������� �"2�ae���?Fr0�Mg��:���@K_c�-���x���1�+���>�Y��x���a��R�<��(��>�r!I�������R�m۶i*K 1];�S�z`�A�8�#-!��3�A�I .΅�"hp4"�q��=;|�ˎ��0������~c�|�JAǂ{��+��_E�S���0��c:b�V��1SN>��|rKs%Բ�'A��ۅ��Gsa���u��$S��Q,c��(�o{ �ɺ���������.d�kR�J�&�* <�W֬]�+I�T�Y�e:�N��6Lą����49� �7�t���J;���I�6H2��x�
���l٢yG ���q�NpEf5`�ܑ���p��\ԈfYKm�93�p��Y	��[��V� �0���A�i,�<l�
��C�j�bH���D;ܘ:�h�ΔL��4�������������c�DQ��	q�r�~s�a�<��%�Mo�\آ�7r�,\��;��cTǅ�1��;'�oN��%>�N�dOl6S����8]KN�SsS]-)���i��?����SH"�#X"�Ѩ�#F놲|����4�Zo2.JW�����SU�Q�*�
(/ѿO�e���Zo����X���C������?�����,�d����N�����Brx 0���&�s�� �6lP����5XU�"bsu�	��Hb��T�qR7)QT2�pT<8��Wi�`��������Y�eX,bڡ�x�k_����.���j쏥������yC��]� �u��cB��P�z�pH^�j��?�fy�:y�O}Ɯ�,����D��G�AlݺE6�y�a�k�I;&���-n��<$���+�V��ɌVӕqN�Ľ��%*��W�xq¼�H��O~_��H�
�C���[eϋ(1�0��eX�[��+��qҭ \m�һd���i�݋�a�~l�TO��o�,U���~�µW�8V�� �}�k�����`mJ/�㔪P|�����Pc �.��'f0�0���Pc�҈��l�����0G]
���|��s���8�%?�D�
���ZY"q�h�0ox���V۲ap 0J]#y�\����Z�!�g��i�J�u+��f�������xg,1�אѡR*�Jo���3f@�W�W`:o�T���?W����]2<tD
�b��j�>��P���XW�f0P3?����f9n�9�d�n	��9X��K����s�>��7� _� H�նo�A3���yC|y����Γf貔���19|��3�ʥ���A�b��.��K.Q�
5�����Z����K�@LLw�xu�ʀQPa��ΦƤ�b;�(�3�_y�zl\�#S�� �h�'�ö׋��nh|�%	�	�7Ζl8[gB�da>�.t=hVN@ðq�/����P��-oy��p�z��䤑M�n�lT��E���n�]�xܑ/<CN[{�T�jR�c�2&=�>	¢�A��w���$g8����^��hr9�%��#��NH�qQft��.��Z��J�]��ǂ�<Os^pS}p¾]g���s���]ق��Aw�]�Y��5	#�T��_��������37](=}+e���%�sE��Di��D����*���7�Q���p�
��&�^�O�N&f�>q k�@�Ŵ  vu���0��ׅ���،�f|��ya��R�to81�
����v^0g;���1�`���K����R��
2b�ep����s}���	�~pTc@lc�Y��KSy2:,���o�CG�w\w�|��~P���Uw�-[P��S0��]m�!�/j`�����5�r�I��(@�����c���5'����QvfLD��ᩤ	�%��6��d��~>��d��Ȁe;�f�
	WW���b�D(�Ұ�;�U�����|�w�I^}�:�$n���:2��1B�';T����'� ��xF��o|C3�x���cB�L��+-���4�j3^���s�9G���.�/񼸨n�q%3љW.xիe�V���͢��Au ��2�=�VFZ=q�`�X*@O�

�y�# �����1��� �=�EB�C��&�r�3v�z�/ˮÆ�#׾��r�Ƴ�H�\�=�R�%����*�&�M7��?�>�cϑ��X�~!��Z�Ɯ���L�)�SK�|��3��ɖ�4�C����$66PR��(�hE��|*��'�#C��� ��������o���$\Q���B�%m�F�9X�|�f��gT�|vK"F}0� ���C���j�ꆁ�Z dۥUki���QË��0 j+ �m�]gc����0�#D��GG�sww�,�]jf?T.}	����&�B#��J�̐K6&����� U4uv��^`� o4�u�E)(��`QEóL	�aG�Ql�j�բ�9G]�
�ɞ���W�R(��q�v�0`s^YC>���F(�rA�"��Ss��2�R3$���F��o�'ʼ�� ���V�?��@��/��� I��]� \N�1*���֌����<E=�4�����_)Fz��PS�����N8r�5o��V����~����2��GU`�����) _���f׈㱁'�_i�L��k�E�8p>X�~�NJ4��ڌ4�m������zG@�~\r<m$���u��S�݆	�c��ƺ񼯶���C���vyp��1C�AXN��6=�e�#H�9n���`��=�Z <���F��$U���h���իW�c��_UU\x��rҼÚ3*'��4��1���m��ҩ>�^I��7�Y��̘�4OE��(�N_+�����^Q���,�*�d���:>��
⌗%S�5�A'�|4��+��B��?���`��ַ�>���W�E��:^ ,Vʬ����	3���������ň�^���o�G�Ŏ�B�2Ci��P�HB�CC�T�uȆP��#�^�3o������6"�p\g^,;`�c��g��n���m�Ш,�d�-f�p�GI�RW�}Ǖr��uf�#f�n$���<z9�!mCL.���%�񔵬BC[OOY�v��r�]�I�5�4&�=��i�3#`�
�&|V*�R5P����w�m��,�l4H���"�5l�>�� p�+b�R�����a�TI���+gd��{�n�u;Y7�0xtl�f�p�+�&�rF����l���0�lR�,�	І \�6��a	�G����+2�z-��5E�Y��=��i�z�5[^�.Eؾo�R�a)[�H,訙�r}o./s�mFiƒV$B.�J�,�l�X>�W!�����w�������a�:�I�/pF{���p��+u ߫��Zə���L��u�8�]��.�i{Eثvb�]�3��ZT�;n��av��f�d�t�޽gwa&r��s��!60c����KVb��	t>X�}��j��1z�3�ZSt9a�8�l0�x���L��k�&kVwK�ё�ډF���U��w�j v��\rɅv��h]B��a��H&���W�z�&9p�jƴ!l^��ƀk�*X@�c�Ft�}Y-dpI�� �|���U�7���M]/�����`a%�&��z`K�P�.��L��8�N^!6�0c�ho���%/�̉�����C�>�3o�G6k3P���8#��f�t	ܴ��Q��.�@����/�J�;�S�>h�d�Ri�hJV7��Oh�=/Ԥ�1�kʂ0��D��U�ȴk�I.��,6���!���c0�oɀǲk�a�f|�1y(�+A\��K�Ы9�%�&Ԣ�H8dU�v?�3�~��o���b#F(1�0���hP&�5p�2���`/�ʳ�C�'T�����̰�l�A��۱=NB�"�v��.v��e���
ɰb�e8�<�����m	�m�C�d�� t�p��<%�����;��N?��׿��e$62�����3�f�.�8�!��;����Zal��e��r���xE�D����9�����$���1|ė={�����ʿ��0@\It�KVʅ��L6l�,�jA��T��	�1�`E�m�ZWo+�(`��#�ZU�(�*#�@����/�O�Se� k����A= �
B�0�wbڝ�{L�>�1��X�Cg����Q丵�/�Ӥ=H���i7|�Sdͩ����v�B������22[l�9TS4
|�q��)�/lU�*h�x@sV����W=0ddT�R�����k*g7;zNϡ�2�z���{�,)���dd�%ʽ[oאK�)�z�Itù��r��a�a�xH8f:8jخY����1g�UW��zVv�8"Q �.Þ_H��bdT��.��	CM� � 緼�M�w�K1��f`�ƍ��g�����4M.��{�,@*D�­1��< )	&���`b���1���]
ޭ�֧%S�@�q���5�46<�����Q�W���iz>���'b�`���@��D�!��@��Q n���xȀ��׽N�?�|M������w�yg�˂�Y>L>�l_G�(P��Ǝ�&~�	{w�'G[��I%Yg����r��bѩH���c#����#��`��}��zV��L`G�B�a��ˠ��/�\1*	�{�W0䫮z�zI ����؏!�XM�}�ٺ��k�y��3]Ѩ"a� �
j�B�rg$�Ŗ�����W���a&�)Kr��ae�o��W4�-"�1h0�0���m�f��@( �3�T���x���q,Ap|���~�#�aψ£��A6��j�v������M1�tH��}�谖zA� ��A��9 ~�J��\��j"����� "߬$R,��f�r�[����%W	Md ��{����1z��3�Q<A���J� �
 @�E�[F�# �XK��X���Z�� j�0#Ѓ j�'Ӌ�4�[�*�xܡ��ry��u�}����I�q�K��0U�/]>(��|��iш�1��64*��P�c{�xA�ш�1�ne���́m�5�|���Z��m�{��#���Tmd\JT'C��K_#KJ����J�����{�O?�9��iL�	�{G�KS�	M���e=����͐�-j�� h�#�[jcCK�s�Ӵ�fm>�I�'���'O�'*K0h؞zz���茡� ��ؙiob p� `#	��h̳�d��c�j,�+o�\R0��EѬ�x��	 CK�(A&qs7�x����4�%t/�@4
@I��x��2�)l6����l��m�+N���ַ�_��_u6�;�� �i����m<���MA�v�5]��W֟�/���R�nؿ����zc�lT���@��K./S�ll1jۙղ?"�#��ϕ��/5�-�Zݗ�%�dhDd�Hu����%Mx�[(��N�8�˞k@ژl�bF�Q��>�W��W�{���El!#F�3�[L� !�*$�O`â������r�2%������)���Z��n����Q�)4 �?�p�P5п��@���ҵ��I�[�:�K�3-S�Q���I�c��M�����5������w�*�x�2��WF��(��1;ʄ
��
"�\�B*�]�t9R�*pT<�R��0��g��R.��z�e��f�4��Be<	�e��Z��|�{���!���R�� G��2P��f5�[n�E-��#�T����nE"��(��W�?2d�A[S��xއD�Rr���& L�\�ׅՑمpcL���7�$P%@����K�.�m�&�=C������N�n�mG�	������n����\�����~�=I�;�&Œ+a�O?�t;izG���\���}�q��D����O��/ɑ��a���/�B)$KZ����a��1�RK���$�$\d��![�1o�!h� �Pi[X/��+j�t�������F���4@8����Փ��F��t�F��(�=�ܣ���p�`��t�t�̺q���g�Zb�b�v���
�\��������O�o�2y�������T^Օr���Q��� ���AF8�2�`¹�R��x��Ы:�P��ȑ1�η(O?�O�9o��
��QU�Y�J	p��G�3)����%I��	!���{�fDw�$�D�	�� -A�o&i��JX�]԰-s���m��(��t�����#L����F�����Ibv�#��IC'�r&�a�N�v @B�wG�@;����'& 3���3�����y[���;�1�Z=���4T���!����3��G���p��cN+�%�s���(��
�� %@HT߈Q�H��=���o�A�8��B�*w�X-�4��G�=�EŜ[�h����e&ۡ'�"@�`l7��x��A�q��-�o��D���t��'�5�ˊ��VR�l$	��P�	�	�V;C~z��4�����!�M'^����%S^��G�=�xiE�$e+�:Z�\���hM��ukd��^��	�F2+k�'4:��xE�"���\G��	-�M����)yAM���a)���c>{�OFd����_��F1��;�D��h�U�H�^I��m�I��u,��b�h<���`��,��[ u�+�x;���ΤF�i��m~�#�:,ms7�RLg���Sh=���Ͳ�6�O�lp���.�ț��Z9}�Js�5e�����ۼVPȓF��rѺt,����%cY�r���(w�����0���+H���t����a�Q�
ؖV�7������*�e���k8���m�4 ��m����i'������
Ϳy�������W_$�>_F���oH�kn�%%Y�AA]��¹��2]7K��g����Uv|�����V�%�Ε�����=�<%�m0+��`<�KO�Ig�
�)h�iE�:I�l�j�6���,�-��`ʻmwޅ`��9����Y���r�\w�I{���kd`�82:�G�{��F@Å�HZ��UU��Ē�ͽ$ryy�L�B��s�(��q�h.n��W�s��^s� w�X���a�}�[8����
3�b!d*�k�UO�U��pڗ�H@p�}@a���YҨ��&���hp4/tɮ���ޗ�S��}���+�'}��_;��b�X�#inkʼs���*���o�`�R���3$�>�TʮV$�`��nCnP��W�zz*j�����X,5UIƴ��I:n���$��L��|�$l��C���eɁ&U�hؤ/?���Q� ��G�J��%w��7f����J϶ *�\r9f��T��������/_�Ï"��z�R����.����H�>f��"�_xN0G�1\ՌN�Jq>e:㺵Js���)��Ubs�l!@��jvA>Ɔ#���5�����ȣ�J����+���74K�����D',	�p'�c8�8'¹��2�N؝��Xj���Q��P��[��CU9rpL#��9u�iV�������Q-�nV��Ɛ�m ��u[U���e��j'��Pf���L8.��G=��[�k�B��;�=�Tn.s]6W�G��U���=*cպ��`44ܐr�Wg�(4������)��șq./_It��JQr�a�%�u�ZS��4�;�P� v����n� �u;�-��خ��v�9[��h�ߵ��>w�I��LY�PD��$�,l$��+4��&J�-�I��pa���Q&L�l�윞�R��J����2:��˨��<�s2u��C��X�A����eI��3�_�¥c�Xv��oZ�dfq��S��d�K�z	Cfs.����
^B�ό���O�r14���{��J�Ud����s�շ��a�F�s&c�d)C�u�L�Ê��b�[&�aUb k�� ˀ.������z킟�1�EG�d��$���a��1{zz�Z}̀n =�.xhHZϭ�՜�ņFBR�(~G�
�Ff8�^D
��l��j�T;п��!8/R�m۶��}�X͆-� �cr�%�ȩ+��/c�vH
^Yv??,���#AL�k'�aU�\���[�	���<(x���m���_s����(�����JWπ����@���$w�nB����Gi����d���$��l Z�s3�Ta�c��8����-xEl���W���6�+�0�u��o1��3a���&��PNA�4\���(�(�2�#�rc�b�ID�����d(�<�c,�^���L��kց�I}���=��v�{v��Y�j�,]f�����e���X�W�è���!륯p���2�U\�9Qn�w͊�e��+e��k��2#��,�{�"8�l� �w<I�kV���s�	��I�ƒ��E6��DJ\֤c}8V� p�եy�H��w(���cH��c��"��� =/����$?�b'���E;˄����:�:�r����~
h�,�����9���N�c�[�7��;��s�g����Td3_;��L�3����s;>,6 ��m��dQ1�����|�;?�姊\y�y�Uꑣ���<ui�m�M������Aƽ%�s��\���
�7 ����i��C>b��3r�+6��ҵZ�hp`�2������Wj��昧j�Ł��^�n���oЂ�x������T�A�3���F�!���r�RG^x���e�&� �ׯ_/7n�ԙO<��w�}
�L��4���0���.��eH?WR����ޛ[z����Y�K�}E��,�UHB�Y�&���ej��$q2���d<N��$�q9�	�+�8,�)��n��lV�f�EK��u���Ϲ����{���,��=}�{��Y����w�+��x1�����ԧ>�0av:���ݽ�,(=̗]��{�2�=I�u�<��:9��9dÂ2�d�����`�u	|F��]�I������ҭ�}N�շ�b�W�SZ �����56PE-�k<L�n?ŭ����LZ<:H�ƽ����|��7��[���q3����t�g���n:vl13�L�23^�2��U�y[�l��:�x�С��]Ď
̴w����Jԃ	�b��|!��`1��Lވ=���ݟ��g�b�A���1�y��:��p�ȌwRQC�; ���W_�����%5��vJ�U/� Tt `L�|�/{���������Ed�2Z�������M8�ߙ�]q�tF�s�F��4�ޕn�w)���>�^�ꗦ=yw�͢�5҄�6ƻ^1F��~������=>6���o���{aW�0:rd9}�K��y4��}n:�A��Uu���@�Y�0�5��0w�za ���//�-�+l5�ھ��o-Y}-��|�W8R8C\��XU�n8U�w�W b�
��`Zވ��q��B�TuG��d�3���b�W\�b�B'���Zn�����+��F��1�bԀ#�]�a�9�
�dԏ�D��3ϝ�nF�#��i���Ӓ��V�6G����#���=�Kg��V���r5t�u�J��ԛۮ���%������u�f6"��jf��↶��F����%(������{~nO"���)������!zW�L)���^��������Zv�.Y�^ı�_�����fS�hZ]j�=צ
�R��O}j�'~_�3��ߜ&�\cm�
 .���.�����P`[r^ r��{��ǘ/�݉�s�}hV�P���k�413:">�q��Lci�%[�	O�y`�=x`!�����w�tɥ�(;�m?��T�^�P]5��_i���"��On���V���[�A:ppoY(`��$���bj�T�r����`�a,�{�����׿>�����9sPi~��/�(��z`p@�<N�9F�� �O�g �#<ª��ک�� �:a�Ӛ,hְ�o~�bE���������Y ZU�_��إxO)w/��ӹ7�x�D�s�e��7��嚟��g� V'lֵ뷊� ��j��28�<7;H��ޖ�>��~�^�'P?�:�i�5̬??�p!��$�ο͢S�-K.��1���[�Sth\��}����y4@F?m��ڧz��rQ���vjYԪԹ�"vI��F��4�8��L7-�׿���;��a������j���4�5J����Mb h�8�=I�UJ�ˆ��R�N�Yi��S�?%D���h3��*N~��wx_�)p��7��#��qb�y�0����T�h'l9 �w} :���x4�-�-�8�-��~����78DQ�?�y�+�Cf�!�}�����ɶ�K��H���_������M/y�3�����_�UE��'C�U#�;���m.ޗ^"�lKL��;n�N�h���X�Dd�n������T��g����\��Y?�T5~B��������矕�ߟ��|� EY�̆���I>p�#�-O�w���~����{�-	�N9C�DL?ap�ȹ�Pe�u T�j'�JǞ]�I |�q�� VQ��j�Ӣ��6[#
����J�{��Ep����=g � K�U��P������b{�7�]��r]�Q�����¹0���������ƸX�^�i*��p9��k^�Ͻ7ʹ3+~�<8{R#��=��H�J"�VI�<U���$b��[d��h=K44r���T�	&��]<z�ȸ������v�"������n�yN6Rg���؎��/��@3-.U���>Et�ra����*��!w�|�+�}�J	 }��^W�v�3k�H���Z*�b<� ��wU1�.�<&�%�h���[ �ƹ  �����������[�R���� ޣ> ���}���RA���*2�XE���y���<�$��KGsM ��y��P:��a7b `ٺ�hԏ/zD�VTX�,��XZ^z ���I���X������{�M�Z�8o ���/"ب(&��bM��m�yy.&o6'�);�`����[�IVϹ�eO�ux�=�N�� &��4���L����a/}�ۇ
�Y\^���@"�e�f�\�>V�N��M|u-Q���i<#����+��+��ha� 3��,�b�DW�6d�u�yX�ϫ�W4*y�5br0>7�x%�Vq���ye�~{�l��t�ܗ!|�H�´���d\��bu=�N����C��DM!0�.���v$�Gv籜���ă����u_��O�E:�A��]�b�L>W�@{�(r$��%Q� %jy��K�V��ʸ����E]�j�0T5�*��=M5����I����C��Oг�Qi��Y�}���p��jYXN]j�5g�����@��}��<�������ԧ��g��IOf���	�B��B� ��x	s� >��a����// Ѹ��_��_M��dòZ�$K�i���un�cP��u�߰^ū`��5��'-�@�a#:%G�ca����]E}���g�C���9�������i����.�@�f�
��`��ǃ�q�tǝG������ئR@+���#�	��E��䩨� ����ϝ%��z������"Fa�EdZ���u�ұa��i�}��Q��jUE�#n�ކ��M���`���@:� �Ġ����N_���Ro8�v��W���Z�J��5�m٩�8!�vQ?j8CB�s��$aF�I81V!��=���ʈ�bU�-%�9SU��t�[2a���1��;�t�X��JS��aEݬ��q���*������s?�sE����u����I7L��9 !�z���q�U�5h��ǎ.�ߙ�T(�D,/̏4d�͉��N5U'�!�
�'篛�����T9�хq� 6�kâ�@A����n��i���zl5W�ˣ�l:�o���}�53�f��i��+u{��U%s0 ���s}����%����__t�	� ^��/�B���K_��d=�*+s�|1߃8��*=u2�zL�w����T	�����fba~��0&x��߰LK ���/ܴ"1/:��A;Oe9a�Oy�Sʵ�h�r8\�{BC�=G����c�V���y9;w_a���ZNS��}[IeY�n35ơ��;�!a߸Kc������x={_3<�Z���?��	�vr!��>��p;�&s��0�ۿ�_��0��]��G{i���+���t�y&\������'�u-�p�*6a�Q?|�_,ċ(]���[��������19�	Ŕ4M,溚V�^���o�h͆���j��R�#3wX����������V�\X�5�!��%�_��&��:��"2��`��À�d�X75��XIaȷ�r�:�4�2p:�n�����b��G�s�:����k�]�9������/�M:t?.xc_�̊[�,�dq�2�<=����L�i����y��18�tD#��_c��Q� QU$kv����Ltth�5.zi�&��w��=�L��6S���XF�@���a�xhu���UWѥ��t���$}������w6��ką��&k"\7�֫�G����R[�w�1|ٙ��xo��g��y��c
� �|��a<�V~W��.~���RZ��I׿�����D������kj_:t�r���嵚�d!���R&;�ɜ0��}��������da�>D�џ����xЪ���b�c."	j�S"�?d̮9��\�:΃m��a��i��= �k�
h?��9�Fg�ܕO(:��sh����u��Iv��`���>|���$�G'� �)�n�p��x��_]������c_����{
�}֞�g�{ݖ��]�Ϧ�G�������q�S&:��V)-]�p|��8X�N& �7T��G����*0���,��~LT�i��B�A}����P�'i�L�{=>TU�QF�`��p�İ�hP@���gU/���	N����9�*MP�|���Q�V/��-���;�s��ϣ���B6E���e���ܳ)5����s�-H��<����@#�qv�H��;3Y�휛n�클w��|?���᠚�s��
��b_��hyȚ}e�-9�����8��:"��+[UltWaɟ����٫S�
��0r�1���c��K�诺�:b0(;(*�Fw5��3������Lam_��m���{'l��N+�M�/
 �VIgG�'�k��==' ��Qrq���:�I�Ȼ���=�%�N/}�uU&���|�_|�+�
�K�V�\���aqY��|���	�eE���=�š�Ɂ|�^���|�P�[6����~ٲ#:c�����S�]�)�9�ދL32Q�aLQ�u����q�J��#�T�yd�V_�Y�z�D�d?:�K.<w��7,A<J~e�5ת��kՃ�di� ��IdA?�d�3Οh�	� �5�'��1�W��x�H��習���;��u^c��kj!�3c��0����qǹޜ�(j4�o<�)
xUn.���д��է}�[[,%%�$��F����cc�N��a\H��^͋��΢��b�˼�E�/��n�_��0��.�@B�I�p.�n�ݜs�M硎` `����?��q�9�~��	 ��3�w��?������w|/���ki�����x�̍˸���p�*�{@�G�υ(D?�@�L��������6�}d�ѵOp��h��Ah�4Y�b~+7(��5Cb���	�Q�$0{?.n��D�n����5Q̶��'?���JUo�%���M�׍ȹ%<�����_�ӯ.��q������� nbq#s�� 7A��im�0[4r���Gy�U�����O}6����p��x�cӹ�<�����d����_�&m>_�SЇ��<�����@U'@�o�1@���ߙ�V���{^�_ԅ`��h�h�9U�bK��r��
��Ro�Q����93]����	(?���"�
]���O �u��7�u�v�s�5��l&9�'���an�=�9E���6l�Gü Wf�L�t�Э�ܜ^��Wd����n��(�bW-3qq���l4� �lP�0h2w�v�;��0�3گ�GH�=/}���t#�n8NP�;>cK�^9�qa�Ff�y��
�W��2�"G�vL;% �G��q�,�MH��8u�)����5"��ܜ<FՖ��(mE�瀯h0�*/��>c�37P����p^���OfU$l���Yn�;����,U�;��̀��S��?���L���� �H�3{��oHވ̀��Zq�g&ܠI"�wr6��C�;�L i.�p��Z�7S�!�W�}�1�Ҝ(�ɑFh4�K�Q���Ǆ�����ԙ�&ʰ�ȳ�FH�������9(�n4��X����R����\�1H�΄��Q���
 �~���0,7B��$N�i�w�f�4�.��QZY��zG��G�^���Q	Ψ�q%jn���ˮ����7�'�('��G?g�&��)�9�A
pH �}��|0�H�'Rt��.:���rl�L6&㤟�`6���`4�����S}�s�0>��0|��F7�� �|�����I�B��'HMH��ؐd�qSQ�%{�) C@���Z.���/�'j07�>ᚑ�sN�ec^k�+�����=��}�	r��n��e%�Fȋg�3���X���^��X��T��d���֓m�R�;@������R�mi~�=Q!��.�t����VW�\�j7��h�q#a���H+lB?#�b��ߌɾ�O$k )�1`��r3�|�K�.k�����i���=��	�pY��qb��Z$7��}�U?_��xy��ޛӏ��C'`���V^���O��ѿ��22u�V\U��.�-�.5���#�o��]�1?��47ߩvw\�y@�����]|K��Z�Zd�47��X#��%�3��cq�|8�`��=��b���5�y=@�	���sr=�'��1n&61�}��pO^܇@��`� ��K��T�6�,����*�(F��l�8�RB,�8��3D��碿8 ���>�*��d!r� Td��C�ٍ����FgF=;cʼ�xv��k�q�A�����Z��@|]��+7����^釾aL7�i����y���u�hlr|��V\c�H�ֵh�%�0������-_�tZ^9��W�TV�Ro��O%-�Š2�>��������L�N���$b�c�}�ܠ����\��܏���S棛�7��������4���Ä�P{ǖ]v,B��8=3��;@�A1؉�Z���� 8<��� L�2��������X��L�]�RGk�ĐBrZL�ѱt���k_���o?U<�٬�y�\|���xK����c��+�s��Y 0A<;;����d�y�(3��Ȩ��::`�o�0��bԡ�W'Ɏ�(e�dt�������E��Z�z ��4��� � '9�x�\�  	�`��Y����8��XO�7��H�ȸ7�ɴ� ��/�ʋq�1�[�+�2^�J�^\����Fk�Uf)���z�2q>4�,�v���M�f�,}�Z�J����l&|��������D���jc�(���u���^���7�Iǎ�*n��3.4Y�_cCl��h�`�C�����9��l|�w���*PؠKQ�<2n�ĺ��2/�|�Ӏ���uPI4OGe|�h\�����a��Cgk}&�{x ��i@Y���q~ݓ\�.VZd/��5�e�F �<��n�X�巼8]x������4���.�;+7"sX��D#���a��g�0� ��A �=@�Ŀyo Qt�t�@�
:��d<����u�q�0q����@�_���7@������)++��α�ȸ��m��c��
��: 'ǨnBtw�	�	�@̧Ap]�	аy���>�=�T��{�ч,n���o,Z��A
r�`�m�9�
�G�c��&2�ڜ�{��$����w6#E�`4P�M��J-�M���dW��#1���m��7��1F7S	W��O�Of��
4�:�t��OM���_������ݗ�^N�),���3�ɿM�յD8�$9Gy�����$��x�zt���s�����%��8�W�	c�ԤD�9"f�~��eW9�v���'��ڤ1�&�L��Jv��]}��.R��04���N� �N�\����H��ufK3��dYJGg �<#�kp0�1u�<��[�d��hX1����So̱.>����j� ñ���KF��FR-� � E�n:>���cf�WU-<L1\�~���Y ���L AF
�D77�Q��T8��D��F]8��Y@�X� �̒��&�Qm{���g�"�2H��	�P��Fù ^���D#z谈�
��G>�w>3/�~���s��K編 G�����������@�7� :�W��Fǎg	e����=��I��{Rz�eOI��q8�%(� ���u3��z�5{�@jڏ<���{�n*V��Q�F��-~�M�괂���r�Y_E�����;���71Z���X��7ͤ�c�<yVґ{o/,xi�P�`wםKiϮ����V��-�T|�["�.�BTsL��04&��� ��,� Xu���H��Tt�R'U^[�'���ٟq�k��ا �WG���ʱ��\�c`|����s��Z�Z�#(��k��Gi�DyY$ �U34[=�Ϡ�@����ʽ�QﮇC]�eC%�􍢪9@3�2 $�����k���`7�=)��F�8+��-�:D7P6DI���0�w��\^s3�3qٗ�{9}�����9���RI����!=���46SoP�0X�������h�٪m���X����<Y�:U���	��E��J���^w�W���xF7��4�I􈀙�K���.>�.��|��t�m��UG�u��ؗ~x0FB5*�Y�k�=K]Ɩ����+�5	\,,,�	���{f� \FE7����䥩/s#�ݱ��q�����
U�?�������q������ת\x&�	��S]��e�����P�%����iaG��Ёj(� #�� r#]Ԝ���mi����2���ߨO���@�uݬ K%#��|����W\1�ce�@�õ5������_�}���;679U{���k�ԯ3sԞ��J?����P�;�+���l6ͥ��=�Oyj:�����-�O�Ae������Q�3��~��\��8Y�\��hC�<R���g#p>m�9��6��Uҝֺ]*�������؅, ;�X��3Gv��r�{���ߕ��⢴�'k���8�5>n̂U��kTV��+�0W�A+J+*��M[ɱ,,U�|����vk���;�"��C���T�D��!@ �y�� 2T��H�� J�h��J0�����Q�j?*N�o��c`��b� �1�9�}��9@��M��{�e�</��Xm����,un���x��Ϸ�0��o�v�zэ���=R��� ��g>c��yO�rO܃���+����mie�xu3��ՙKwޅ��0�u�iiq%s�,��D��_M_��;���O��*�Oou9u�k�ݴUD����<��u+6IQ}�D�9n�_�P����V�Ś_��q*t�悎�Q[�f��j�	�R�ޏ��Z9���n�ñ��ư��2���x���ΕdR2��;�LD����H���}I��E	u��'lN ���Ɇ]��O5@�0Ѓ{U���q�����p��waEi)�J�� ��|n�7i�.�2{p֪���N���e���Pk �|&+���>��g}J�����oA�<ԧs�z�"�s���_�{g1���G~ �㬑Q��:�is�TZYi�@�k2��H��k�lg>=p�p�x�ymeIs�f����q뭩H�7S�P��dY��{^/�;&1�cں;�6<�>�j���CٱQ�w�����hQt�܈��)z��]���w�?�>��v���ۊM���͋t�'}����ˮT��UڞQ�r��\@,���F��K�]��_�{ݗ�C������{�u��g��M��GР}m#�	���c�e�@�H��]XV� �Ȟ�q�Y�C�X]4��n�V���F���7���]m6*���ٜ 4@��ͣ
�ee��*[�?���+vC�9�q�T��=��<�c�}Y�����97� �q����g��8�\�f��'�u��%B�7���AZ�k璟ɛ,��a�V&��iqeX<%�>;o��"�s
��5Ɖ��/nt�s�"^�}�@=��u����I�N��Vmk�Q�7�r6��Q_Y7Z�p�e�N��q���Rv\�?J�P��ꫯH�w5��0ͤo�ݽ����+--c��)���l1QRe�{���X,�7%I&&��hp�K�j�c�O �jl
?�:���M�P�F+�6Lӭ�H"��d�|�ƌV�D�@8q,L̠��	ȹ��Y�d���� 2���Or��{�J�O�HI��
2Ґ��q�:�ܜCC����;�99��bf�������a����>�zƠ�յN��^.1/�sϡ��q/2f����y��o����d2��F�w͑�}%�⫟�^�����\� ����F8+�uj��ހM4K���q�8#Q�g��W���؅A��&���}��(���	��)u� <�'Yv�F{,���+���޴U֣�L�"���Ț�nRu?��8��1�W]�_WV�r4O�t�y{Sp$�u���{:s�U�fv��"Q����Y�k��i��gq#�i��j
<7� zpO�v}!c�W�u��b�w@s��Ⓟ�j&Q�xt��h����LQ>NJ~g�f܀��70<�w��ƨ�t��i�y(�4�Ѧ��c���{NXolO�1X$����iج�5��|��i�IT�9��3�a�ul�;��^ �^ݸ.���q�D��g��v �����!Qo���XIg�1����J����=���'�o#ϫQZ<�(�`��crS��~�n�]�~oJy��<�u��@c�*?U��,�����.�{��%Ap�E}��w�G3�^�1 �{����w;��0���F���#��ZlG���zb�]`u�v���2>]��M�ڠ����{��(�w�Bz��.K�����Ky?�J�'��+k F���*߽U
Q@@0S��ϲ�Q<e�I-�ɈQ�b�f�p���Km����n@5`�-�u"�J}��o�i�z�&���N�E°�wu�����7cqu2�9N��bۮ�9��4:�ˢ�k}�5��G�l�C�ޓ��M�����Q�yZ��G��j*��T���&��������:P�p�W�e��m�=��m'&x���.^Y��6�����:��e n5�A�hI=�və��	�Չg&"y�v��w�F~;�,��h�(6hx�^W?΍�]Ռ�O�G�VW�Lo��^�~��^��ҽk�;R��0��󰪶<����/���K.�l4�ϚU�{dN���k����0����������2�4���߭�[\ [o���������A���e�ݴ�nv���u�'�L��5�	�H���l��¥�L#��|�ӟO��ޑ��I���/K�?[ x~>��X&@�����	�/�wd���h<��� �$��c����mc�e/��ؤ�9�!"��6a�m�j��G��(�ɮG���&vH��d���F����n����=��\tx2>E�1�ц�H��L��ٕ�{)}�c�~��ǧ'�����xHL���y. b���,�Z*�4����]��x��x�C쿸����"����xYr<W��~Rډ��F`u� 6��nv���Zu�����F`_�~��6z��4��U�l���0?��>����wI��L�=�?;�R�#HPe%]7Қ7Ud���X���J�UPۊFN�EI3�����|����͙m��{)�C;:�̄��l��`[c ��y��C?5�;{�7 �X�aS�?�u�և�
02߭�u=My�0a/�N���O1�x�:`AM��s�Y��W�����7�M�K�4�!�CO?Uي�ͱKZ0Ѝ6WG��U��F�G���
S毕�}���$�ƈ��KM}q���!=���=��6E��g������`i[�ش{8Q�?۩0�킿�4ͮm#��4��ζaq�Dm7$��Q��������3/�n�B'Kγ��[J=Ԙ���iϢ���\�+�*��Y�u�F��f�+mp����_�fTc��*��k�������;�AC�`X�,�kT)�V�Ki�W�^v٣J�E:�/���N�E��� UQ�&G1�.j�26_�-:����Ź0��c��q�������/3%z����G������´ɜ?����Y�ze�h�Imb�
�e�5XV�R��s�S�z��'��rpC�Z����^@W���&�h��3��a\��Qo�O�O�}n����|�����j����`l#��Fg;s�e�o�JDe��(DXE��BԯJ���8�1C�����׾�����>������+��h�ǥi��P�{R�^y啅0�1u�\��� 1 O�KL�Ͷ�)��v�QF�E��2��	a#�ݳ7=�Q�MO�3&��`������N��YB�2�X�Ɇ�\w׏�����p�&U6�bt E�?��?.�jb��Xbm��ĿF�'$�����^���s�={h�~�2̥����ƨh�[�[���L9W���`�L��4�Q|�( ��	}<�~�
���a�s�2���I�Eo�6���7hlv���Է��&��9��t�����O���uY**J2�eN���ۓ^�/H_���gr��slD�Ƽ�g;%0jee)���KC�;���\M!��iQ�F<��,�ɍsL�)��X$h� `�qx�@H��v}qM�#�]?�9�)XCRx�m�JH�`?�ߝa�@�/���xEz�S���@y���9���� X-���z�K^���O�tRa"zV��Dڋ����u�1���Ό���>s��6�K_��t�����yr,��ե�UP�F�P��p\�5�b��DSfu�F����/����
���e�B�-�4�<�����RLS�._�z����'Y'|*m+�jlu={�|#�矦���s3�]7����a�Zy�o�
O)~���	 �ٵ��qՕ�w~���S��t�E�j�H���
��t�+(e�x�i�z^�a��3�� � f�j�pǊ�G`��W_]��
�`m��|J����{)X��1�馛
��}�Cw�v<bn4LFX�O�9�I���?���%q�s#hS`f{� D ��l=���� =P9�ܮ����{�yt ��}(}���ۍ���"U\�z[o�\�B+U���׾"���t����y�V˥�܈���A���H��	Z�6
;��U-T��GU�F#�9$��琨_/�b&�k`�zf8���g|��i-�F��'�m�з���TJh�����ot��x7A�I����rNKKi����[�>��\� �c��ֆ�N&����Go־m�b�#�Sy��J�:�=�;_gO:Vr��t��/J^zA����b�[]=���K3}���� $����Ӌ_��w�[5@H{�;�1I�dȼM&R3�������;L�B���"zd���/6�I����a¨#���w�V������Q��С��y9D=�D���H90����t�;m I����e/+�!₺S���O˥���;jW:���F���oݖ�;wEs9�J��]�����g�9i���q��x��/c��z��������\��j��J`�d�%�ƅVw@����~ְQ��,t��ͲNG;ϣD�{��xZT��bܘ�<Z������77b�"@G�����M����F�q�|��p7������~��<W���=i���]EW<U��� mU������ �?��?+��@L�Ԙ�Ԡ$��T �%8
�dyf ؠ���գ��z��������Q�vm��M��N�Ǔd�ߪr��t����
Ӣ�0�J���������≘��c�w$���~��������=�yew2��:��ӛ�[Â��i3��a7����O~$?ǝ%yLw8 Bno:t7eY�dqk0f�c�`������B/��Xj��b���gdr�䜗�nu�1Z��_f ����l+]������~�3ݝ�h�L��T<�@�b���h���+螥Ǐ�o:��^O�Y�:k�N�
M+�d ޕ�����#�#7|*�������ƹ��O�:�y�i8GC��6�A�^%g�)"�+�>��t�7��X<;����s^I� /�����D�Dc��zt����<��#���O~r���k�{O�O:�7;��Ǐ-�7LG`y��7h�.ߣ��0�$�7�	�����s��a� UX3����ԸP�b��Dy@x�A׻2�=^,��A��[�,�lwW2J�;��z�H}���Dp��P`����cSP����CYYd\����v�m3C�N<{=�JF�/:���M4_O:�]��Cg�9�c��=��!�y����������yMt2���Ez�kϧ#�g"p��^�x����Sk�R����Өt��3aUeJܣ{Я�گ��O�_�ksx󖷼� ����rN}�G�R���g�:��F���H�@`�C�Q�BBQÊ5����L8��Q<�IfЏ8�s���&�Ao�>���6���` ��P(>��3���ท���e��X:�����{�{Kgt�����N���
�u�U&%9�3C�Q�O�!��!ї�ۣ[3�g�|Ƥ=��~q��|�I�j\b����g����1��� ���!?
��V����P��7^s'�7b�H���S������77�9,Xi�;+�u�Y��$N�y]G���:uuDQ���Y:�f�^�ղ4��n����i���k���-@�_���&x�j'�cLpϽ��o,j�c��g?��x~>ӥR�˹�_�
�f�i���4�D۔BL���&�W��6�U`o��`�F�?Z�,�,����������l�UԈ�~3���b����`h��\Oy�Sҫ^��I'�[���N��z���]��a�:"N���]>�Z��,n�K/���ӘOݕ=yw�?�g��#�
�� <J�zz��|��؜@$]��ͤ#�� �A�z�gN����t��$�}:��MR	.����3]'Y3,~2���5ZCD��l�w�D��Ѩ|�����M�fb�����Yo�Uo+uB�Ľu����8s�T��hB��L������g_���\,7�T��1�s� \E��<��5�����t�5�U ����T��?Xm�g׌^��4�=&��:JVR�n|f�cQ\pW��Q�qj	�OHQn�^1�IRv�V��Wr�iD���b�[��s�P�3hQ�Q �'bɯ�ꯦ����(:|����g�z���4�M��bzы�Lg�����-�fs>�����?�'�:��j��W���/� �Q�$�9�>���V#�d'Ϧ��	�,�v\h�?��Û�u�T�
�N��9��֯����1���T�*Rm��Ҁ C�a����H�G������P��������4��/`��be�8���h�jN��ʀ`����tn^Co���^��g��YI�n�v�����l����h��Kq��\�'�nhu�6���/#���3D�����e���7}�zrܢ�>������Q���4�
�muO�7�n�5���kV7�5��wח{l5��x�~Y�zN�ĺsˢ-?��w���\LX6L�-�V��!�b[£R%�9���ܩ��E�Jn�NZZλgcWIFR"{FvY;m���m����lOQQߡ��1�}�p�~����QT���
F�i���ТԶ]��@�o:����o@�o��
�3E�����ck &��1��s��� l�k���y�?�Ò
��ꗴ���R^G)�;�.�i��N^_�y"W�(�����̩0�q�Z��(<Pi�ˢ+�U]1�`8��e�GOu��F�K����@�3:H�� {su��5[�Q���7^̣�I�JG�@FQY@�n$��Id�E�b8���Aa��/�忤�����x���S�{&y�@�p�}?梒�w��]��G�N����R��Z,�s�3%�)Y�ƽQ�xF̬yKl�Ec@l��R��4&N�i��?��(��F ���F��,+&������i�#��?kL[7)�)���[�g�f-���5%	2$��9��"o�����N�� ;�y]3���X�Ъ�Gp�B4�q[��sh��(#&��
 f�*"r�~i43�����8�7�?��R1p3�G�/�/��/n�b���/K�ܝJ5���KH�s���&8a��qݲ����o-�qG�x/j�4��{��__6�?��?�����T��E�UF����Q�i~��I
c����j;�;ɶ�N��7��(�����e��1��y[/*���w��99�w�R6|f�Z	�X�%��������b7gpaLl|S p;_fASE�:f�i��n��_�n�t����%O&&��4d�..h�qhGs��;�����@�Im��;����X0GНi0�`L޽��آH����4 ���z���UND'�[V7o�7~�� s���Q���4bT�_nhQ�S/���@$g=p�qtKs���G�ܕj��J$�)�����.[\<�n��O���7~/����ї]����/���5���R�s��� �e�;�=�)��ozӛ���jbw�"}�Ā4ab*�[G�n-� �Smj$�����)u���	�����/Y�mt����,���=�:���ݭ���CE�a8L���U��������d춵�����L���|�L����7_K��c�׿4�y�A:T�s�@����}I<2S�Χ��f�+Y�e�yY�GЍ%�l���nH��F]�|i,D3ũ��1(�D[�}Ǘ�C_ɜ��1Y
I7Js@ˤ�}�g� ��Cp�XT�1�Y�}1�Y�OՄ*9ƈ�8/�G?�u׵���GԵI�3���CZ�d"���f5}�7�C���y��M�3Ӡ�7�h&1�RH����Z��d������Dʰ"9}������whх�y	Vq<R�D�9+fG��͚��`�5�8�n���΃0MŽ�ą���yl��{�7?H5QxX�G��N.2` �cd,�6>�*���]�c���g��GL$�	��\�>TvI]�bL��ހR~7K���G��_ �LY��~j���=UG�\�1~h�QO�99�������E ��u׶�g����bFOU�=����dT�O�G�����kxV}���KSt�~������y�K�[�$bb�� �R�����ѕ������
*B4���'Ԋg�Lj6f��Z���������轻:�\�2��ۈ����^��i�Ա�y�$ B����}��.}�Z�_�7X1�d�a���9�:s3f���/Y���4c^���q����Ou[;��F�q
���L���z��x�v����M�f��e�WUh�-�����>P���y!�DL�/|�El��8���7��t�'?����L X1zb<30�=:\g��:��,���`�i���iq)�`��=�@z�c&�gH�s�ʢ�f�Ԩ^��S��2���/�7�c
O�l1'(!��[��\� @K�����o3��6ꍚ��µ`�0.�1� �p�_4�>M���`��nP��Ju�lWM�l�����cY�(�l��Ak@��Nj7��L;R��	/��#.97}盇��b8"'L��Ȼ��>�id���ɧ\�Vz��_����� ,� ��9zaT�GT���i�/ǰ�+��`!T��4�G��	hƏ1��p!؅���0��lХ|��0��۱�^�w��~���(a�;��$#�����N!β禠��1�����fq��Pο��o.�9���hX7���-�F�6;�L�\z0��%�N]�_� ��f�z���{q*蘆zrv������C�YZ�1a�VRIo]�L�aEU�V�a"�D}��1M*c���<��s�n����-O��'���p\�HP��{�~ ^��^�xCf`�J��LMu�L�>�m��舭��� ��֔���r"�=��g=�n)Rz��l+�3��O/~�u��dl�I�|�h�
o��TI�k�Kq�:F��G��!�}��^{m��AU�O}j�p]]:}��Ma$�%�C�s^/��'�8@��%�N.���oi��#(�93����ц<��?���{�t�ŗ,�?�V�Šk8q"3	���X;����Iq�1�,nM6��mq�G>�ѓΨ&{�zhL�ed�X�|����W����ͦ��}LZ\>�fڳi�t�T%ܝ<�*#\�3��2�*6�g�[�%��1b�A
&2��&d�ɞNT'�zz<������T"����d��O�C ��������@4VG/S G�!�Vw�aql6�}�dqN��kV��5�� vӆ�T�ek��Z���'y��3�`�V��g\�Ĵ�ey}��3�<���#ŧ�����������I}���-0��V�@y���EE2��&�s���֞����#5���������;�#�ӯ~�u�6�p�����Ύ��^&�jeG����z��/|I�ǗIȎc�"��.8DU����ތ���G>RحF#�TY���/:����4YX��D���v�)-�.����%鬳�(�t[���N+˽<A��Օ�0����үQ��l?���80F2��W�i��f-�" �;��/-���)���ۉ�~�w ��5�(��<�����/��,Y/�!kG]vd�����l ��p�
�	�d�l��j<g-r �=�����:hʹR�C����l/��XI{����v��鑏if�r55;Y:Y��n���k��j��ꪸi�o#j�L����!pT��y��5���y�hxv�XHϸ�2.�	}��a�V�Q�~F�ÆŹq��5�Z�C#�X=��L�֘DUU~�3c�gb�`w�ywȆ���*�� �b#���_�bQn�� ���7t3�~���L8���Q�Ϣ6魎E�n-�����ay.e��a��׿����oڃ<1��مt��y@gw�!���n���+nzD�u�U���PoV���{��aA0A�ie�Q|*�������7��9�\�C"�N7�	�>��O;���w��2F���	b/�k�˭���K��3�p`�Jr���Ƴ���1�[/^f��.9�˔�fb��X��E������' X&AA�eʅ�f�`6[���0K����3�%U�#�����|��Ԟٗ��=P�� -�ߝV{˕zb�Ve<��^!46|�� I�6!0�������4�K�����
!Τ�%�i)CCntd\�_^0p���w�l�������k���qI�CU��7*��X����0꾜:��a�kW�zе���"��q����%ȸ���E����X7���a$ ��濺1���Ci~���*��O���Jlj�˱�i��Rߣ�����Eo@Ft=�FٝhηXbD㿑��N]�y"��^Ի�7���=�O�`gp���@���FBc-���%`	%����u��ArU�l�w�u�T��F:�z;�t�x���D��{����Ꙇ�� �p0�ڙ�\���ff| ��MeW� �������6`�N��7���FĜ���&��aM:��T�5�$�[p ��CUi��O��ԙ��E��������9O8d�\�v!>�3���[&��&�| Ev�<t��%�D��u���ۛ�PT�3 �;��z��q��p4�}�����O��9��Q��=�A9��ü�������
�x�\ԑ]2	g���Dܮ��j$���cܙsQ�|:Z]']7ј�z�0�!"V��l��74�&4#�8�u�� ����%��M窚EI����>��-�G�>��^cl:Yg��]ψ��TUmW{���3��Ŵrt��9X���_��-��/s�V�L$'$���� ����-�;�o6s@���(�<1(E�� �IA)Ƅ<��qyŠ��n�Q�9��G'L�j⍳菂�����swpM�nn��6�T����h�h�����u:��	�P��j\D��������i%���l��#�9��V�$q�lU��A�\1�������4`����i1
�D|��jaEN�4�o4���K��<�Ws1_�����orQ}�C�S�+�3ݫT���<��=�C��=!y��6##�p5�O����I&4�yu���J��ʌuZy]f������R�]��vJ�!g����J#��-���'�U��>T�#TI��FP�n�5͋F_�hߊs=[O�m�;���h��n��\��ϢU���-.$���4�n�.78�fLL;�D��5T�pK�/��u��,B��H���^�5O�cu�-�5n���n�R�c)���?=�nէ���P���;�
�űӛ�;�ft���m��H4�,Vw2��vԅ��Z�Z���)��1��(�,��*{N^��#���6d���F��:��sˈ���gh�����k�K�]rNڳ{��Cbڝ=xg�Ӯ�*�{�y�T�k��g.�������ّ��b���t;�y%�?ٱ��J�FqN���ʃ��{�T6���|�M1MuSh��	��`T�6֘Ҵ���\����J,�W�u}�h��u���&������G���E=\��h)=��'��g��r�;��sF��H���?�n�-R@��xs��19�9#d�Nds}hMvb���vYpl^C� ��wJ�q"��!���4ؔ4~q_|f�\��F�ׄ��t�ENc� . -���2Gn[ �ngQ]ǵP��ր	��@aY�(��&6��uy%��e���=���k�s�{u�(ޞٓV��t<3�]{2;���\���SXtņGE_K~�z0�FW�W��r�(J]p���TM���)��,�.�Ӣ�'��t�@����Iw�N�G}��wu�R���Y@]����ˤ�R���kO���0H� &���Iˋ���=,�<)�ͦ��F:|��#��w��f���VTaT��R�A���ޢ+�(7MdU��i��3T4�L;��]���玢*M 0o�^9,t�$��F��u�ܵx'`��ݤ?S�ZA�y��#�ٺ!a��/�fߨ������G�5�]��/�^�)kp�Vj��_����)�0����J:��FqUC3�j�O�+�t������L�=���cX���5�)��Q�ZR�8���������M�c��c%xu�1�6�Y���{-7��MAx��M��z�3�)n_щ^qJ�(]�Q�'{|/��3���Ȥ�P;�	��J�k�K��>��򦏦K/۟���G���۝Ť����®�<��lK������i�I�PWO�uc���i��Ӫ	�Of(�>O�q�~u���z2p|�ȯޅp����`�F��o����� �!�%�3_>l�	U!���u��X�����6"�h��k����:Y*kfiq)}��_I����ӓ���t��Jǎf��ٕ�-��(����-^��Z}�~ҝ/�O�F�C�_�?�Ҳ�$V�u7ʺ5F;�T����n�:����RS��-��Y�hQ�R���5�s�~~~�e�^;2��ǧ���Z�TϏ�i������t���7қ���~�.�g�yR�������Faヰ	�~$���|V7C�� ��d4ҝ����`@k��D���TtC�'{O�5"��m�2��$ǉ���A��n"��`%�B\;4Y6�|��*�~�<�$̣!��;TlH0������'kl2y�`�:��bجW���g��+�7������}��ON睷7u��|;����'�Z�*׮䫞s$�����9�;��ű��N�w���:j�5rwJ�~S���(ߘ\b|�k�_q�h���q�(Fx�'��,������_��1�zu�s)�=�O�<I�����&=�W��>��%���2�Gg|���Q��x4���N8Z��i��t�<W��  f���������<��w���Qw͹�zy-�g�C��Z�ܒD���Moð���)F� �sN��P�{�X�ي��:eذ�]"Q����Xj�Y9���Ψ$jG�<r�h���8�Z��v/��V�3ж��LN�G��z)j'��>C�=U<��umu�`���D����'8�q<tџ4�Tf|0;!VM��1�Zd�3{��^p��:u��|b�M�RUy��,�u[閿�3-/Qv&�R�S�=Wr#�$��I��Q��Pn����H����.q'T�m;�[�,شE��N�s�r�df7u��j9ݩ`�օ�� f���� ��c����9A��djzr�⼀7��]Y-/Z]=8MT��o�RN=zdt2;˼��b��Iw�u_&7�t�E�|+�ػoWQS�
��-k��N�7Zw�mbE�k�q�k�uf<V7��)��MA��sv�dQ�ڼM��`"�	±	�u����ؚ�q�E����w�-�r����R��f暙)�"��ԙ���"���3,Lx<l�ᜰ��u?tq4�E��rӌ��p;-2���9��4�Lk�C-�պ�wBg��׼�ll]r�����a���	C����bXSg�a�k�� �a�a�oX��Du��wDɡ�`�@%�kZ�����Un�Ʒ�$ٮ�g��m G@���5O��y-�:?(�H�Cz�fk��+�̠1>�f4u��ApZ��>#�����ql$�Q]�mLQ��e4K���l�gQ��-�.*�xg����c���n}���3�����T�k��,#���3��52��}/�ڛ!x���K�����t���ґ��y�P�1�q�[o���w{�b��v� W�nd�Vգ�h\U]��X�!l�EU�j2ϭ�D\n(�\#�ȑ`a[+`����9 W�lh.�h����P{L�8+��p�>�&��I�F?�Ra�|+��g�s�>�wϥ�_��t�p73�R�����JZ��`<[�ёw�0��cp��r3 ���g7��X#1���љQ��wx*lxsn������	�t�2Y�����|ŉT_Q\����Z�U�#G����]�RG��ܮaz�k_�.�p&]��+������r�s#ZM�/�r�4O�S,)��������� �e�i5Ĵ{��	6�	ڨqO���QԮ���4���zO�> K�Q}Q�����OY����wo�(Po�$K�?�b �k�G���f���Ͽ�{_I�����������lvP���ٚ�l�\��4���>����>'}�w����URY���-��J.��z����]�˳ҷ�	�9��a�
�p=.^�q���MAx8h�0��0�:�x1)�Ư��x���6M�+�C�k���D.ӌtu ���E�;�^��̦��ܚ�7�^8�Ծ�$*q2ڗ�7TK�>��|�l������C��h]7L�	]d�&Y����4釶���ʄy�f���}�<��l�uт.�#ޏs��PQIX)C�<���Vu�=�#�9�I/%}���h�,}1�2&6[5���n����O��s��tB>_|zgJƲ�\�����ݕ����Һ���:�J��]y�<��oN���E���$��.}�O2��\�`x�x��޴K�an&�(�`7�N��5"EG��O���/�[��t�f�0���AT"��٠l����h^O|��5�\S�g�'�(͝�&��*<͐T����~�+_O���L�+���);�K�~����6*�\)�R�yTÛ�M&,�g��o������IFK���͌s�xND�y"M/1�Ĭ��ɫb"��PĔ�Y������`�(���d7&׻�K�{%F��K�ϴ�i3���6�^&+�O��̂WZyø'}�K�ʠ|����p.�ʹ�{��t��invO��-���8^��h;����������I�Y���s2���<�a�)�S��-t�Pr�.+!���j�<��^z��W��{Τ�9�2LE+�3������:M7�tS9>:��>c�����/y�����t�UW����-��9d����o/;M�B��}|�����A���[I����Z��Z,9���y"��Nǎ؄��@�DZ�Vs.�0e��P���x�p�er4� A��^�<�����9����Lr��i3�>��O;6��Ģ�3�+ L_@4��i�\� g�,��E�K��G03�}��v��Jȵ�t����B��R�'
Õ��c�(j�Z	�ڿ!`��"ޗ�8�_��{���tÇ>��A��I�wq��OJ��|)������)��:I�d���70���^���� %%�ԛ;M�M	��4�~��+��#8w�7g k0��G�Z�CI$��<-�Q{�h5[�����)�1��,�'�ܓӳ�y]ڳg_��ٱa�N&��x �EN:�T��V�K��V]�j��ԔBd�?���.ߛX<V��X�1od���|�]��d�{h�Ҿ����f�f`����nx46$4�9XmuD�iup3�D�&��n'\��O�\UCXN����t�M�T�V@��  ,N6ve��*ki{uۀ  ���+nz�����Zt�����PE=�6K�����Ozz0��O�ռn��u�Z�MGC��s��u[fó��S�Y�UW�K�Kl-�{�/fD�oc�SQ9V��&�8S\�����7JV�x�3������k�9&����=8l�l����+�O5 ƚ��5��d�A�6>���yIf�ץ����j�h;1L@����`�щTL%3�ᛑ-��#�9���`>N\��h� �3�peۃt�H��bR^L��2��8��9�x$�#L�1�-7�J�<`�n����n�r�	
�7bB%��E)�%�j�ZQL��+{�0����^��Έ�6a���(�\�����8ǔ���0������?��-",�Ρ8m��lR�W=��'���[�HEs��H�����3N��B'��%��WRZ.��о�v�=#8X�a/-����[�y���+éj'��-�K���������x�;J?�[���CC�M�o�q�4jL@L"�9�U�P�tp~3F`�VQ8�͕�v��d���i �����~#?��t�W���~=���3�;Zyo��I�P��s��-�Z!��>�/y�K�w��Ǽ�u�+���b'�X��0�z�	�$�LN�����GfJ�~��-<����S+l���TJ�4LH
>�A8�t���I�	u�y�K�9D{栬PF㦿�0M�\��y^�E����cX��0�EC4��ҏ��wu�y�GI��晽v�H�k�Ɏ$��௚�r_���V�r$]x����F�T����.ܥ��<&u����/�{������ )�fc�!K;}�ӟ.����P3��1�>�&��� 5�;*��1:ڊ"��g�������1c���}n2��N���h0��/�,t�W����)`�t*`�e��{'+��Э��2QM�����:)asF�=�O}�:Jv�v�Xz��H���I���4�����ݝ���/�Gjj�	��!J�V���|����{؉T3>��殺���et��Ǩ�nX�fF���h�Z 0aĬ�]�ۚW���7K�RSVE7W��Ut�C��)1'�a��sG76��Dl��Z	�5�܉��s��RF�f�iv�\z�/�<����N��^1|�;s��qX�\j7����uG+�_���n�ES�B5�A�1}�я~��R� ��RmK�q��� ��
��>�s�^�(fx���3
 �G�h���X%qzK����R��L������!|��a1 vI� 8�BG;���� ��yk��s�k�oD������_ˠ����[�^L�������<@�i+���{�&��K���RvTJ��Gm ����H �0�y� �9����3�h,66]Æc����s�噙��!��t�YG�M��:\�M~���]�Q"�𞱁]z,��F!H�w��r�2��N����]��^<v��/9��~B�������L:v,K2�nI�ngf��R��y��ݔ&�rm��7 Q�#ρ�FX�)��4�0�h3�����
=�/��➼4�2���ê�X��;τ�VAv��^p�y�#��~XtK�nR<�)�5�#D�B=1��,s>����ꜛE�e���zX)_��W���J�]�1@#����X1��=������\zFz�k^�f��<p�8_��I�L�s��@nϰ���EO��&[cc>���U%�x3���0K�u?�m���h�tB�l��>�����@+; s�z��u#d�3���"F®)��ҪM�T��y�7��Bj5��K��0�/9��I��,5馛>�>�gQ��ЏN�3����?���l�uE!b��}G��׿��E%A?��.�U</�y�w��]�>%%<�x�3 �/�P�Mi���Ҷ��8��q�]C(��
Z��q�y�s�����bqgh��}��W�� ��Ibuc��T��xH�-����B���qC{�k_[vA���t��t�;���"��qq���2�.��#�/��>������;����oo-�r���L�1�e���"��DܿO��Qׇ���ԍ�X��X����I�J�,�t=&;�`�Sl�ޢ��{B�C2�'��em1��x����~�1�&M���;�K�X�a��fܞ��z��L��+����=���_~�3����ҡ�{�7��t��{K��fs6���R�3>-����y0ȿ�e/+��.��oxCynt�|nE��!�XHb�b1(��(�sn�EyN�Gm�=�G������ڈ���UG4Z�ҵ�[%x����$���ۀ�$oc-��;��+�1������"�y�~����������芟��g��e�q������¤�sh����ӝ?�7}�O�:��U�K�>��H�b�+j�F����Uʲ�Fy�7i�Ֆ�"��XMs�[��m*)���&���b�N���&�Ci�~ΓY�^G�k�s�qm� '�I£
�{9���K��;2��
�3�%�Xa���`�,q}��XŢ=Eo	����õ$@T�"�a�;��owf�sdm��U�������t�������aw�u�T�f��3c�W�,�	(�̪��G�e��������˛���"��;�,+��������x	YS��O�~�����S��k�2H4�L���8����'=��PG�G�V���ʺ]6]���k�ݍ��S��dwٲ�_d
ՀV:a:#�C��ab���\^ӿ�ɕ돆ie9�C?�/��<IF��[�H�_p^>���� =��\�u�-���+�? � �Rg�?���.̦?�fA�U��L��۽׺��k1_�/�L#�� ���h��4�kØ�7���r�fk~Ƞ�E�,��^�}��Q�,[Vա�� A��D�M�!l��WW��J�b���]E���݇Ұ?���ޔe�|��������\e������7� �w�H�آ�J@����'��5�)nk "�D��^�)�|3zOhP��^��	)1���UQJ�4Wv���R�hT��/4\cavRw�f-��."ѰJv삈I5h�υb�c_�җ�����I7�pC�\X0j
\G���?���"]�y�oa~&���H�>��tɥ���fz��}�J���+m�����yo�F�>�g�����:ӭn� .8�n@�ewd0��E&b��9�ew;´�[��
���Pώ�z�-��c�y�v�q|�<,�A��xǄT�SC��W~�p���O�_r@iD_�6Qݻ�s��\u��<R�k�Է'23l�Rg��.zę閯ݟ�C��WJD*�#7e�Z�̂���~��9�x�$���7��<�9�?���T�A�~���wxWi�:q7>]cـb��8~q����X�X���W̭���l�s;��h��y��r*f�|��z����;o�ܰ��sx�)ylԁY"����������$5y5l�I��|�3�)��23Fm	LS��ưL�QZI������_|Af�g�W�+CIU�QXq����vU�S@$~�ӞA&<���T��fM���YwK�Qb�m̱���T�a���*�#�ى��F�I ]�̀  �� @��)1���[�.�c��!��ڊ��kK�aT�`��QEp?H�lJ��j����!�W���if���ϥW����;ߺ?9�/u纽ci�ފU.-/�
+V9\��+V;���'�X՗����o�v�P�oHƀ��싸�}x=n4���x*�4�����}�mu�E�b�*�&/v��@͙�+
Ɇe���Z����g1�E�gXA�F��D�<�'�����u�G}w���)�Y<������t�#���_qQ&�t�b�U���**��J/�~�f��6��D�u�0�L�M�)����n\��N�im��4����U�O��{���(��J��!q|��z�H}.�D�DI�s�o�g���Q��X-id��2�<n�[��/�a�f�XmF�6F���C� ) 0��	k*��}�������e�|.�������͡�OOzʣҿ������Ng�ufa�Ԥ�u�a�_ȼ��p�IG�z^?~�����/�R�PF5>plԑ��Dn��TS���Iċ��Qu�����d�����}#3��p0� ��A����shb�b�1�4�ޱS�!�L�Cǘ�'2X�75�:6un����uT�E��;*�|~�0]}���}�.���X��Υ���i��?-�3#u����q���6N�=c��:˵�.�N����f�Fu��'{�h�ޮ:��D�`��+�v����國sW�<@�8�0b�)`k�M��vp���ͺ@#ܭ`aVW�	���_e���fL�!�s��@o[�_T����iFs��������˳s�t�Ż�Y�^�n���L�qSg&ϙ6*�n��y-���R��0�=��O��C�����Pb��sLc���8�Ք�ԙ�;��6��&��W���y�Z��E�q@����m���F�v���0��i/z����+�t���ID7�>Fk����/f�ѱ��7����Y��q7�9\��E� ��� δ���}���T�$:gG�����A������-}�;�����M3s��޻���eί���/����ԊZ��@�iQ���+����K{�n4.x\`������������4p����:�Ό��.m���ν�U_��A2�Q��	��L�f#�dmH� ����Ju����m.c��8,�kFC]TM߀6b���y��3��D��k^߼��t�_|=�gKY�Ngwcj8��Rf/--Ri��:YR����fSM�S�+=����ځ8��~d�yғ�Tp�M�d`�Ȍ���Ȳ������r�ʪR��$��Ҋ�B 	#$�	!�1k;lf�D���3቙��n�{"�1�&�=xŋڣ��2b�X�&�RH�U�de���߹����n��r�L$���Ro��9��?��1�DԲ�1A��zL��Jrw-�asc��T��v4�[et��)1,�D`�+�ޢ�۽`�{��Ŏ�������Wy����L@���F�dI(�tg��}��Q�#����
�ӟ�L{��L��¿�@�8��}���h����/3w�Y;rx�*���E�;��7��Zb�]���s��(5����yc�6!��� ��Vmh���ă�V�B�K o.���}��7v]S�y,iF��3G�$(.��LR��浤DU�`�(E*�6��������w��W���wJ����pkAj\�}���K����LP���-��_ ����	ϡ���ȋI��趕3Yx@pUL�����?�~#��/�R��ؐ��y�5�p#E���g�
0��_G�)���ø"���F�cUdֻ&�u�N��N�2<�Z��؅0������;Pc��i�3qxϮ)[�De�(�D&U��N�k!�q=�0�J��@�
��#��2����[>��:'¦�C�?��V �r��ӧ���O�f�`�Y�\	s\����K��f�5�d�^?�@=HϹ�+��_�^��u�RE��T��4��ȧ�	ӭy�C��km(\
D=��m��@�����,��Ԥ����"� #n?��|�"���"�6�÷��.���3sԢ�N;�jVo��|���frpWm���|�*�}aN�D{K7���+�^��\W�\��j#a�������g��0b66��J��ؾ�D<�P������g��+:��W�͠7���8���ګ#"��$fg���ِ�'�z)B��'í�!�K���L�Ag��@���X�M^I/X��r7RzLO���&� �$@��85�OڲU�jV_���#ǭ:1c�V�z��v��@�2�IA��D��p�C�\�QQ���8J<��_K��:��ꈥ����leD�����d�S��S��B��Q�{��ET/���6�ݻ0-#� ��}bڎ?a����rXS��%o�	��'S(�j��i�c���*:��a�b~��T?ZK��BlvHҤ��qc�C��y\�{�H��s �T���O�6�|<W=��
�ЩY60�sQ��N��k,��(ّ�XE~u�
t�F3�`���X�Y]�^�Ʌ���|gO�-'v"j���:�!��e/pK�u�7K�L��'���UJa'���!ڝ��}�f6��Õ�9;���?��#�:\m>E �6��>J_��+�����J��L�Z3^�/0՟���|//-��x� ��Bja�.�>�l�Y8%��|���eo?�n��%v���5�#z� �Y�I�)
@'P� v#��<Y�|`�����/��{�Tr�
9 U(2�-!0|�Y
���RܗvQU��<P�XC����W֨v�$�^���I{:�r���ZqY1B"Z��>�������_�'q��\�zΐ��@�K���޲\B޻ m��@����]��a�hu欓�;x�����_{o��ɤƦ0�[Mc}�,:h5$jM$����������a����К�R	m ���rΫ�._�����z��h��>�e܉�O[��`�j�6o�loy�+�U��>��k3��T�@��Y��rS~r�z+%�2f��e��sA���u��l��7�
����=@����x�8"��:Nc��2/D�����*�ʟ�&F(��,�m�\o�s�O �Nf��Z�bZN�t�dgR�W����A��%��x�(�׏ϸ��`�Y����Oy�=�'Æ7|��1	b�FY�];��J�c�d�S[�f3�n���[��軒Յ.{#�!Gq1�!|���a!?^�"����(�96h<�~	x�3�j5��rA���m�<k5�X�����42����~K�[l߾zn �t��@_c�&�����20{젚��^T��� �0	���SQ	�U=t�✹&@�Ď�^AJ�i]�������~
�N'�\��70�-��kWzX�ۄd`P#�������yp�� RM����T%x���lI�A��B�n������l�[n�:습���v���WZ��l�&vx5���݇��Q�<?��w��Q4�h��9y��=s�{�]��=AF%��ǺQJ��0�[aݶ�6Q��q�ngE�x����W��]q�Kl�maΕ�L� uv[�Z.j>�G��(�P̛����9W�DEo�(F[ ���q�W�e,S�>����6Y�`/�&]7l���p����jt����A��~/ZD�����-��	<|��>�Ĉa�P�E�����}Z���[��'�x���w�զ'7[�r4�6�<l9��WJE� M4���\�0���?�/��V<�sL�gi�Ӧx*�ޜ�?�Mb9 X��d{3"�z��A��Bs{�d�)��v5��i�����J��r����ޯ��/�gs���_�2H��1�p30s��Mo��n����&)�3!^U�DEb"���H/=��5ߕU���1�:����=��/�^�#!�ƒ�-2�Ҟx���GK��r>�8A�*�����Jr����b`� �{
�}���&s<�[�m[w�S=i��������ο��p�J�̇�N���CE.�G�y#���'�7��P1<�/B����s��h��o�ɴ�EYW�zf�(�X ���"������e2es-�]T��̘� `��>��v`���n='���/b��S]R6�����^۽߭�Z�&5�"D闯�&WL�_ᑷ5q�2���^Hܸ���=�y�s7�k�.U�>މ7��jJ$�7�sG~��8�;�{=�����Hw�c*��E]�o�~ǿ�ı�yX2e�����_&I5`������ӵ~ވ�j��J���@9��I��z�i�������$�C1��O�q��j�<W/	�or�7�&��U��B/���@�Y�7h�o��"�� .h�X�_t_������'҂�����W�)�iX��\fv�ZSv]�*Q�011�3X��^hԛ��Oe* �YX��ʞ�d��_�
@��4wG1"а�?����������=��Q9Y�U1��I~2�z�Bq-���������/��}8퉙8�ʕ�.��۹k{xo��t��V�~}9��"�<�]�[�=��O~qkg����{ ��{Bxg-t/�d��-N�a�i?a�!Ë�:��j)��_ۻ�s�ħ�/�G?���`T�t���W1^��g染�,λ#zfE��v����E���Q7�'a��}�;��Fy��/8���^��:1��j�
�����[�;�EXj�+���Qs�8��ڄ<���or�I����,pdE.�����Z�IEU������{&�ũ=}�i;}�6{�O���\p���(���u%�ig�o���2�[��" V[��P��s�꓀ƃ��"�i<}ٖa��Un�=��Kaq��f��C�ߨ��B��p����"��9�9�^>�gy��1}���W�U{�$��o vo��QHs�?{?��}nkKX�[1,���6��6��j?��[��~hG�խ�:fI�a�f%��$�eU����W��=ޟ7L�YOZ�\�߰�S��r�=jw�R�k��5�c�up�����;��sv�%[�y/8;L��(&MLe��-���p�J��(2���U\�9��yqT���X/���_��׵�3�F3��},r��V5>BI�F��g
�;/m	��o��R'���6z�H/�K��P ��`��I��W�����"�΢$�LR��jiZ�� '� 5�L���y��߿~������y{Ίf�y�! �i� ���)�Zq�x�f�r�.5Ǉm��1�QHcA��rF2��-�P�IQ��5���S�m�z?Q�����v�i��~��sΌ9�X�[���U�����Y;v4tvi,	�X����٢�������@�"Ǩ1й�ĮS�D�g���^>ۛ^���{q3� z^-N�Q.I�|tm���;���{�aݛ�DG������˟�!xc�f��]	g��� u�R�)SB��n\/�2��Пٖ ƍ�V�{ٕvڶ���ө9J�g#�q�,J��d�5���Z\�K6���AK�?�v���%#�hʸc��R��*Z�}���P���z}�?����そ-�,J��a�}�DԋA�*ۉO�7��7�f�UȎ��r|M��e'�fƾ=ŅU����1g4+��8*n
zv��w��O��^* q��+��7ho����?k]S����(��{5Ű>�;Iҵ�;IR#�;^}��QR��&�$!���VQa~�VL_����[�,��=��>�����֌I�[��"�N��ju�QNia!l�]���������_��r�Z���.ُt0��r�=��T<]!��NfolO$~�{����b'�J��|������|��B\U�J$C9f��sv`5��Rn�"�S���}<�P�,+��Pa��E����K_����}���A��V䊼�<g\��.W�T_4��,j�{�N.WV*ZI�>
|�a�f�5���>A")r�(ɍ�L�GD��z8��TT�����&�K��J���I4(�����s?r��ү� Ҫ���)t�k���A��aR]�y?Ӫ�����X���i�gp��⮏؇>�ak��Z�bڦ�7�UW���\p�5[��)�5�>�w�D�a�����U��8�Y1LE��4�+�%G +�b�_2y��{Y��QT}�W/����@�pjo���!����ჶ0Oٓ�0qjv����z��l��C��o^I �e�n��D��$�E}��d���s���< �L��b�J�_��m����< �"� P ��r����W���=�^ �$D� ��|~��⺤?����??r�@�������ƈ���8s�~ ��e�+�\� K}�Ky����RO �ܟc g�!<�M�~��D���򒍣����D���&lQ�09U�Ns��	\/Z̪5IY�mZ����=}��0U*fn<ƭ�s�Ԧ�S3n�8R���o� �MP�N��J(]%j��	N8)����pd]O��"�V%d/�	KnT��0�8e���l� Z�<���x�x p#*�B�#�|)}�>H�H�I�3�Q(Iw�1 �<����v�B�bY� �!���$} �'�61�C�u�^K� �~��u���.5цqEu�(Ւ6C�K^���o�̓��92'8_9 ������w�7%�`���"�2/�@"���k"��]f��}+�������L0�h#��h#���+���6����?ǒ��{r,� �	k�{2wi3k��Tƞ́$2 k�q�����_�r{
������w|j4~����uJ��a�F7ϰ�5լ�ZxtSd��j��kA
	��MQ�#KE���'�c"��j�y5�E����E~���}}���>� �+U$�}�+l���)V��><#ի��t��X�u;��p,;==K�3Q�<I�(&��_n�^zi��|k��`�3AI/�����n׿�;"xS��s�+��"r=>�`�Dz@��E/z�IA�J�mǎ�0��m��CN�(�M�O����7��3�ѵ~*˥��W��O�FLyOx=����|_�qC�TE@/�CWCE���g
�3��c����U�u�ߜ�Q�X�w1��1?�r`�q?�x����[����7P����CF=y+(_,m%/�R�z��P�[ 5�q]@S��5�Us���b� �!�2����e�P��,�	��)R�E����l�36���X�h"�&lێ-��+/����\km�=�0��Jo̕��3	��gI��T�����͑�����G�#�LT���K6=*� }�I{���:TL��Vj3~�G��E��讽N�RIڝ�M���'����n��^xQ �kbZ80�k�d�<&���&zB�DDB&c��B�g�g#�������}Q�p�7F �a ��\�EḰ�� <Q��^����D%�Ī��Q%��������3����
���Im��~�?���N�YXԅ�[�i�86J�Q<�$=x��]!�S�aj&�=�L���	�c�Ј�,0/��V��H t�|f����8�9(�8�y�F�25�#��1��X��E*#�a��\-t����VF/Iq�Q���y�C<�r�;�t��}���Q��aé�r���2��܉#�%aOڵ];�����F��/��Z���0��Mx�V�Z�6=#�2�[����I��V�4&��+^�
���ۣ�8�ӗ���1/0e��z��C������|��:,���4���x���Y�<�����v��),a��M�,�Ns�n>�l^t��t��ag:�W�
΀�!�p`�Ʌ�]���j�}�����ʎ��"c����Q��w�i?��?o�''+��u��H�-��h�����ݴ�w�<,���/>m�f��E�jŹ�>�F=p�)���֫5�u�^U�d4!5h����NznΨ�5�����,nE���s�3��� ̢�w�ׇ"�|q&޸��<wDI�f��X�,�é>`�����.d^�^|Fg�x����u��F_�I��SqJ�bh �J��A�h?��E����0�6m� �\�)��?sԵٙ �NV���F�c�[&�3�Zu"H*iۦj����M+U��Z��e`�ݾ;$�P�UkC���������+_���9�o|�#C���I�>��&ȳG�T��넥�{�,��!�0�G ��Z)�px�k�	��(6��M�͛���l�� ؝��yf���	�>ɧ�I�?X{:���.�"���R u�kq>0"����ܱv1_tO�$��7t9G�Өpן��sׄ���l��M��Hy�p�q�y�r"�[=��N��0#����H-�QRzMMl�V�<�Oj�0���a@�O�(�PŰk��7@���b��es�).�k�P9��ec���9ǵ8���5�
��\����yϢ��zp���,\��p�p�������%��}�o='����0�5N~��S�	j4�1Z7m���
���4�ԷT����߶˞s��>繡�%�Q�+�$�����_�U�!�C����s�p�s��%%�o��Jq<c+@FR�馛�3a��5�^�%FI�<�c޾�/������/�g(}�����%��������&���9�X�ͯ?d���ý^�`Lnu��G�k��6.�,nC��{<�������|�#��?��?�7����Ap�StA�`�]����:e��_~�����oٿ��_�߷r���|4ט(���4L� @�B,�|�m�5�G��a<�4P7�:r	[�3�rh�J��\@J�x� ��yϕ�����g�J���E`�$��F��@��a� �Ap�0��o�}��ĸs���}U�$�F	�̱0J 8�7��b��pq\��dh�I�+ΐ�2��8�L*>֟�����$L"�N�n�#�Gn�F����������{���j�˿��&'�m���"��������$�Vyn��u��W��mx����'���}�8Tm�b�Ĥ��c�d^������u��'H�K�bs��{����VXop�k�����Q��������"b�1�i�2�h��XJ�"]��3vFO��f��Q���ɋ�C�̄G��7��w<����"��t�ϖ��M�y�t���#v�'ﵟ|�+���P9n*����fä�M�Vޏ뽎S�n-4�>7,���=�z�azY��E ^Kf8ԟ$�le�l�SD<t��@%zz�"�1�Ƙ,��A�����\��z衞�!b��ay!��l	�7��g�T 9��& * G���Gnm*���K��fA������c��J�����s���稛�Ƶ��n+z�;ٸ;ڱO}�s�������4+'�Y���l�1�5b����?��`l��/��^��WG	��t�a�P�s�=��s57 l �b~@|���֐rxh��yހ�7�7U��P����a�	H�ؑy2LT'�.�{�!��3���#��YF&;��/t�I̎�N�D�a` �{����4zd:����_��x.��E��̊�;>�x�ĂQ(v�DÞzr�]tɥF��VNx2���Rf�[f�r��񐨥�#ø�a���)�P�/��$2�3�@~���R�9 ��� Wɜ�h"j	���3��׼xj�h5�2h�!	�4�>_5s�{���7�q�=��I�r���K�"-|��w|���*�#��!{�|���q��~��:>P�$�>E2�J�)1?6����$fJK����
���u�)�I�կ��??/�O�������8Ό��-�_lzR�ȷXz[ ��Fg�f���o0~y5�X�3|V�E�2w��
a�k�	'�r�M��	�X�t+t�"�GG�k�B)�(�Cް^'H(����u������-�qD8�l�z
0���s�uH���=�)����6�NY)�����n{.:7�T��V�\�ʢ��tn.�D=��* ����`H��wYS;�G��-F���������~�^�Q�;�"�2X�T= �`?�R%� MZ�s�������@T�u����	�5�l�"����B  u��@�W��j-x ѫ���ŤDޯU�О��5�s뙣0��N��ȅ0|[� �i&�����OX'��|c. ��L[XC�6y��ܐ��m���*�:yI<I�P�T$�1��JqTr��v#y��j����ل����J���	C�i���k��хl��YR��N�T4��Kc�2h�J8!������G���:�� j�c��B k�ypF�R+�F��sv؏���p�r����=�U�������D7j{1�b�������yė@g�ܚ���3+�L�mY)yN��?f��kMî9N
�������N�F�v�bëE`�����^y�=���F�4;|�`�/��.���S���0��,��#�/���XI8Tc�(�$oFa��d�+[æ�C}�6�  ��IDAT�{�jS�����ݼ_N8 �8t9���[e�G2����h�XVj-h݂�ᢆn��[o��	_��1�NZ�F,�.�M�Atmj�do����=n�+_p�M̴�Qϸ�Nhnti�p�#R��'��9*m�E�ٝ%���!�sJ�@U . �$V���=j\�3��Î�z����\�z�0�|Q
7�0����n�C"��+i�!\J�����_�cs�;v��^h_r�=��&gg�n"��U��\�U?��i���} �ԋ0(��N~�#�$8�G��! �^]���$n��:FҔ�^��Ͷ·N��ˣ%�m�5�Һ��G�����@ ��7s����� P@����G��N�k�1�<<)=4�HK��\���E�{l.j��]��l�.6�#v����n��a�L����yu��&�KDU�5�"?Y�ּ�B",˫d��s5 ���Z�"�֥���~����b؞
��u�Q��b��:ܵ%|�����a=LN����a������mێ�;�[ϳ�~�` ް��Sf�w�.y��֩�\�ۆХÄ��o��0���>�v�0e��B>�M82�z�(5�����z�a����n�[.-.�xB��&β�A]�:#�_�ThpQ����������K��p��{�[�b����i��{���g��6�t;�|?���|�R;�[��������a��)|��N�D��FgI#l�$@+���Pz?/�+��(�k\��B���*ǩ��Ѩ�4��1~W���{H��c~��+w��p���@�dڴ90@Uk.�b����}���Y����?�J�6���ێ�B��wZRg���|��	k��s< X��{���{��8E4�ە@@�A.i�� o�	�e��Ƒ��K�Nw��5J�v*=G\i���v��¾3ޥH@Z�pQ��nG�uL�k����aN�~Ǻ�կ~5�������Q�|�3���ǃpֿn����_�;v䐕*d|j9|�m9�:s����Ls�\��H(��,�Ч��n\㢉(5�al���Y>�D���E��ն� <
�W�E�jQ�����b.~�/�� U��%e[�_�|�c������8d��MdJ�b7��j��Tmr*��0g۪��/V�2^r3U�� F\$����ߏyq��-�H�X�!�&x�Q_�ˋiz�K�R22ڥ,o���I��n�V��XQy#�h"��:�E����x7o$�3.':ݢ1�Dˑ�G�O�/L�b���3(ɱ�J}PKc�σ�f�-V�$a"a<(��<��Ӯ�a���9g\BU����ë �,�q��ǥ/�q� %#�Oj����J��aTԉS?�>+1>���j�.v9���j��6�g'�B� NNLe��e�I\A��R5��n�gm����|�N�~��̐U�eR^bY�BI�a���d��F+\�X����C���M .�_p��3C�Ǎ���KF���q������{��R��5�Nڕ�#�����p�sϏb�	�%=O��_��1*@C9\��A�NGu�)K��irD̡�G�Agg$���g�:I���V^?]�K�-P�_��j�H�X��Z����J �ސF���ؤ�ܘ�Ae�řӉj�h��o~�+��-�������)�J�s�Ji�Jf�x����(z���&�Fcr`���F e�%Ҙ����T��~������%i7�7�W��>�ASSS�Q#X�w±pɄ����������~�5a�̎���XT��{W@��9C� �|0Hђ��y��-�(�BZ�M<n<55w"�.����H�� ��=ј�n��%�����̎�O1���:��D�d�#a@��1�	���5n+<��ﾻ��ɷ�{pm�����p�u�f�b��J9��ɔ�����M��C�	�K��W�f%��C"���;��+TG��{*r�Ec�8�wW�T[ƵkԹ�8�����h�x=A�_"�&��e��d�sRH�KO�6��8�G�ݳ1�?W+p��#>}�v�/��?�Z�;�
��l�MK���=�	n��{���Ђ?��?s�p�hH�G�-; �8��+�/8�ڒ�?
��:St�sA"������6���^�F�N��ֆ�$�s��2cO�����^���Fu�SO����>���a���� H �`��JN�Ί~"<��?��?�����ꝏ[�|#dD<�8!];&�ڊUx5�r+�؇��]ĕ� �͘O�r-���������~4�C1N~`t���a���n�=[���V �e�6{�Ͻ�~��o��Z �:�Y�&�a}&��%������E����N�5��;�w3�E-b XA�ɢF�@����%&��j'�va��سgO�d�/� |P�����R���3DFGp��Db�i��^-�	�I�XF��$��:���c�Չ^M7���h,�T�'�T�$r�:y�]��^٬C���[b;%NhW�@��A�c٦&7��][�J;2�ɠ�8�<� .��Vb��aI)��6h�����T�42@m۾c��s޶�VH_9���w����o�s�6Mo�)/QS�N�*62N˾��pq� . ���uWK�T�J�$��WG��^�
��ʵ�����w��3�( ��b�b�Pn�bދ��r"�25��dL�sքƱ���_���z��#Gˀ�FB����B
��X�6�T.��蠀����t�ܓ�Jގ�T��+]��q醉�==k؁��ؾ�����fw���љЯ���m�����a�V�Ֆ���O��A�σ��4�ymCkY�q�&����ڷ��d`��
�q]S�sj����/ ��>S� ��T�p�bʊ�%U�����6@ޣ�p/WO��&Q ��6�?���PR�3,�'V	K����Vo.D�����"G���N�)3(
�``v+v!�F�w�*�Ă��ك���׼�78��2@�Oj�z>�ם��Ժ�m�|�}꣟��O�#?x�����ض�;�`i���M�;��,����l���$��X�� �Z���\îҲ�����7��v�������v���ע��4�b�����Ի�*��u�]9R���J��J����� ļ�������B�;`^!��Yد����Ғ �@�)2��-���H�tsp��P\�"�a��v���9%�� H^9�F��
�O�B ���Q^ �{����6��'�x��򃟴׽�v��=-�GIE8�wx���E� ޠ���D�i*�&ʹ���0>��O��s69qF��b�2x��,�� �:�0惫�//@���4�0�!�D;>�I*	�����&�
?1�ΐ�׆��5�R).��h<�Ԋ�^�8.��U;�>3�Ocu �Vɪ���3�C���2(��b�xQl+����������@. UjA�, JVI��g�*z@���R���V���{roVl�����ٌ	���;Q��A���r���ј��Z��o��������c�nٹ�LS�=�q��R|��ԕ+�{H�VjD�2�B��T`�7��W^	~$|.j>s=��Sp�H��ʹ�
�����.��}n�4��>.u@�\NN,�̦�x��b'f���є�V:9�= [t�@� aY�"qB�t\�xK�C�1��AɿP)� �W�|�'�*�z���|Ĭ6�Yi؅�m;N�l�S��ޯ���)��ōN;����ڠ]DE\cYǋM@2 �T%��-v����_�o�*�^�lW��B��^�1[=&/̏-���*F�J���>�X�J �+^�n�a�|ДWcB*X!X�}r��֞NZ�4�#r�t�U�([ϐ7�@�H�G�x7�������XY6�ex|>
��j������O4��w��t������ُ��z��2ʦ���9�T�F�{��h�c��Sk�:t�<�6��r�>����҉k��X*}^4Lx������#�8����+�Sc���}���?�$-?��w\π?6sIMJE꟭o��->E���[|��L_�NJsHY�._��V{�<�k�0��}r%1!�̫V����*�ʡ 	Q^GR���)l]��x`Z��گs��y�c��� ���o���ਕ���ݑ��LD״ޜL��R�+��杘6�&�<��Q�����1�L ��>�s��Џ�;>Y�`�Rߓ���G9����,��8�-�[@��V� ��xw�!4�p�/;a�N���[�KΰK/=�&�Kv���3S5�cXr߻�%����DrX��F�o-7I��W@L�ߚl���&���姩��r��Z#_j��=�H|���r q���ʷ[�ڐ6I?*䟵 �K>Z��_R�(O�����;��RV�%SH�.}cqS���}qU��6IH̊6X�]I�z>>$]�D�/%5��R����7�{����͛lbj2���\w����
{������3b�#\:kթ�����w�����*Z�&T����
q?��m_iE�C�'�(MWǍ�>�����/山��a	b��<�����	9�m��l��Y|�v��������9�7��2CC�'�.�W[.YV[��J��>���X���.U����xx�b��B�X!��6Gq�R'	�]+$T\�mD ��8�︎rp=y���(N�K;j���|�ө��F_�Sz?-lq��bf.�y�bD�U�C��,����$�{��Ӹ*����K�.���a��E��j�/4cy���b��n�풋ϳ�]fss-k�� Y�H���kw���h�h�9��43��+!yRx�P��J��an�9�F��	�;&{�Cn�}����K����&�v2-�QC�������M��i�Z���>:g[gϲ��<1��sP�#N�W� �}�-V��L�,�Sq�J$.S��D@ ��X�ճD��-p����%���(#վw�����H�Tj3��i��y�R�S-7�kN���j���ࢴ8���(Jn}�(4����^��D�}���o�z�r���m0^#�Z�**È��#���FO�jeҞ�7g_{��<�0�l��B7[703��1��Z����3�Tb<����o��Wh� �dFp�˹�l[?�[A��Q;��Z���RWxqP �wT$5�|�.ngs'�W��v�:h� Tu���g�D�F�'7e�"ba�NLa�Df8/���*	)����������1Y<�Q
Pe'�q��	I|g!(���ŕK� (��W�G "}1�䪦"qO�*ݭ6��A{U ק����p=�)�c�VMqഏkpm~�]��~�-\[ܳ'�M`��Xc+���zR�����1��6L���b(�����p�R6�N��@Kܼ�U̢�^�g�ev�;z���߹�����4�Sj�I;|���}���u7��]gY�4��b<Ƣ�/�8�� ��y߼$뙸�H:����\n�9�xUߊ��'��������M���vs�Њ"?f����>wb��'�:Ĩ01�h���	 ^�n���s������	[?��~� 	���cq�X &�^��^�X�8� *�-w 
�)~�J~����$�^zit�Q�@��K!^/������x~���8�w��{"�����M���{|�rJ۩���'ek�$��]ʅ�爣�t�RPEW�� �#��O��v��2(������n�#��$ƕ��MQ�p1�2���H��u�;!���>JGK�i�*�r�+��N�6	t"��"�h3�*T�gGpנ���2^�햔óճ���I�6�FN��X��^I�U��'m ���{yھ��w�G�.xS�Y�ͨ#�:�#q�^�(R�.?�8�w�%^�9�	\�{�����5��sZn��%�T������u\6�S�5�-kwI��-��0��NసVu*��rFT�]�I�"���ʑJ%j���ű�	�Q��N
P�  ����>�� G\v�����ߜOi�����+��"�/`��v���  ~�>�`�� m!3ɺ �.� Ĺ��`M`��T��K{9�� � �r_Tuc�����f��崝1�ܛό# ��*}.?S� ���r-��f��f$� �6����@9�񑏻���w υsy�<��&b�1�;�:���z�$��� @�b�3�����G����9�TX.%�N��2F-�AR�&Y��tлD�J�3ʯz��焇q�ˡnw��	Ot:�ҞRO��*�x�b����E�U{u�#Y�ДA�u�]�n#N���;t`�@����dح��a�΍p�ˢ�?�<�_�D���Ćdܒ�	�L�Z�3�� �D�X�$,\@���x�c��NΉ�R% . ��� h�� `D;��-�K,.�������m��s.`�m�x��q-H�5zv�E�JWʸ�+���u�I;��6p]ڦ�d�4 j���6 `l!�9%cýd�U\3@�̹\������fD{�� ��OWc���<S�XQ(�TO�������`֓�;b�S5k�p�u�<S��;�0*ktӆ�_��g�c�\}����9���uV�R��D_;�	R�TORE%�Ai��ԁ^R�h�@��ƌ�n�B�wB�b*���muc"5���kAIg'qKzE�(�1�<�(~ �u�� H`��`��y\������9'��J%�햛�cS��z��&j%k5J��ɖ���;��G�Y+��="�Mn���W@�� ��{,�0u�҆�Dn?�;:�K�'�����쾺3�	��BC!�ø3�(s@���9�c/�<+�hh�D%��$��Y�� ����/s�Ϝ�=�N� J��xp> H[�tʊ����q�@��sƐ�܇y�J�|T2���U���O�c�#��VF;qb|��*1���޵�����C� 6>�'����G�.���).	s�����ǣv���so�I{�-W��dhC�n��R�[lrb�-,�y&���	c���G%F�A�#	W�S����|�Oگ�. �������9j�C",��]�*�{ch�9�n))U˕�g9 �lpR,�t���*E�%݊&��E���a�8Y����t�,UP�N��]�;`{�O�=I���~�v۱}6֜�v�V�۬�[���1��s�>aϏ&�����A��Ȋ�o�	q�qg�XIO�o�	 �ɨx{�ѽ!D28�y ��3D)U�P2����K[�r�&��ui��^����W�'O�B�űÙ�8SUX��T9^_�O�6-T&������㽌\���r	 �pќ#��r�p>=���4��kr,��o~����I{�'����b#�06����H9O�gq�P!�v]�)��UJ�5�l��	��bpu�[8f�v��O�N�ԯ�����a���\���V�6D��v�|e���@ء�^̋���xx?t�����P�Yv	��}�Oi�������N�'��.��J��KY�Z�U�?��N��w�]�	�B�=��.���jb�kP09`Y�e ����鑊�vSQ����!;��vÍ�И�a�[�Ul~�p���p�eu�'�·*�_�\�
�3�f�͸*��W�B� ~��+_g<�^g��H���4�p,|~c�s�V��3���(��Z�<x�'�����N\���k�����f�zCB\�<+Tq�X��Q &�����9G�>��NT0R�p�Bh[��8��~P�	`�g�ϱ�j,�K����5.�˜��8*�>�y�kȅϯ�����c��-�a�զ�9n�G�m��?f���vɥׄ��u��Zb�z7��"�$ϙ��|7�օ�Ah���}��T\�gc��O�m�k2y6��4/�!K��p%�N�ֺ�r�SI��ݥ��%I2	M��o?=r  �V�5$�*�c�9�ゃ�k����K,�$�L��0&?�0]��2�(Z�����q-���B���"7�o�-a��ڑ�lfS)<�N�QˀXE=#wrP^? �����&���r�J�˱��G8+���� ��=L*��x&;�	�p<�l���\ �de|y��$�ȆH)��\�x�<s 
�gŽ8O�)8y%a�E{T6_ �v�0����617��ע��ƫjJ���C�i�Wp���h<���W�1��1�<��8T�)�8c+uc�x�,�+m�m|��d�L��T%��gB��ӆ!O�u���~��b�l�X�1�O��b�>����w���֨W�~����v��o����R�<���`�~�T@�� ~�y�KV�"���j<4��K��ld|׫M��y��F��#�e�+r��Zµn'�R�s	�!p����v�,����.�k����)�� ��o�ǔ�c�P���cLbb2�$���K�����U��7p����8pЧ?��\^"�(gu�	�,%��v+�;����vϧ?o�yͭ1�O�Ӵ�MC���:�����[��0F,x9������?�X�Ð�X��])�����(%�:��s#LD&(�v ,�ǳи�:
�г���t˼�N�$��㸮T
����C�^q����7��g@�k�l ���o��y1�|/� s��.��`^z��IZ�pO�Oq��2�%�}%Y�_��I��gmb���U�z�}qf��/~�0s�fd/(��u��U�am���S�Q��ԩ/�����=�������T�t+'ӱ��f�oe%�� K�qw�qG�����!)in���{�9I�+{�|đ� o0HA/�S� �1e�W�B���=7I�2@��T�+�%]�*�0���Xc.�i�p�<Q�s��+k\p�E�E���!
�O�!:&�@
7C� 
�]D�4�p��	1F�ǽH�|�7Dq�kHL�V̆��g��'�\�&O- FXDO<f\tVh5�8eN[_�����~�H��s&()��p�^���s�3�OARoh2KO�݅(p�2�
|� 4һ�;���>�d\��(	��) 7��k'5��?�%N^��?�M�`�'����"����K���2
�~�W�\����MB���`L7qc
~Иs��q�0���$$�D!��j=�:O�M�x"�#+��j�yZ�	�0s;AWO4�-# �Fla�y�k_�����7���_��h$��<|$����{���o����iH0���#�y��`n�����ճ�z�W����{G��J���R�8���-���XE�`�����tǄ��Q���&5�V�X<tL�*E�l &�o��oG���^�:���?��k���o�Piw*& )�L��τ�|�.��t�𢳣:��l���"��,�{&9ur��J?��:�/����o4Y']�<Ε�����k  �X%��\�+xC�S�%�{�I4=�-�M%��.�N�~s����w��T	>���@��~kj��W�s}��tw��i�)��kjQ���8E ���&�!�u-�Qu�I94��q�&�st��W�K�K�ubn>����NEIy��;m��h[1x�"�����Q6�'�O�^ �+�XA�"� E��Cf|��К�3���*<�Z�瞽!�k=��Q�^������C�k���@���ђ�p���X�ʅL�ո��K���1=��
~�|�m��tϋ_��o��A;:�����>f��[��.��!#�w+iaxn��p��mb*v����{���Mw�y�i�a�3�r�R��rN*���YC���3����E��G��G�����=�h�c�}"�aM�H=����x�s�
�+�&?�ݑ��Z�i��%�(oȟ�=n�ʵ����@)/���,JUޖ��R�/N,��J�����a�z���^���I�T>�k=�����,X��h�R5��nD�6���U��;��}v�ȂMLZ��C{�S�c�Uצ^���h�;��^��F�����_��CG�J��ɥ�'�B� ���1>��&�ׄ{����o�b����jkN0!�ݩ5vQ�&jUk/�^�'C7s�aW`p����bO��B�iBH��$B�HG�%�R�����ϸ�� ;��� � 2���}�}�*��g`b&kv�ۛ��v�%����1`��Y��8���'^p��][���o�I�*���Ӱ�x�����N�c��ŰW��W��ڤW�J�H,�P`Qz�ܠw��QM��}_�F�߆����v�����1)��u=��k��|��~�-������^m�c��J�i+��9��*���I���DVmrz��Aj��*�5/��~��������q��m�\���P����f>c�Fs`^+i�ThzN��jozӛ"|��}��2.�%T��n$)�5��M	]�ʪ�,TZ��X��<`�6g�Q�̑)�I�_�.jI���S��4b�2A�β#��t
�I<7��g+w��,ƀ1��Yq�pw�}w�0����-G��܀��D�����Rb[wL�� }��۱#�6�y{x0-�7�<��-�Z醋f}*�AkA���5^I�R
LWg��������T'��vع{���?�Ή��'�mj:K�Z)�֤��b�@�D
�6*OT� ����ƜB�yEj�0:+镘6y�h��+�א���_hp�{t|&��C�F6�iH��j/� ��l�F�L�ð�J=Ile�؉����DW��Y�pź�@��)b���$���x8Oj����%DN;6ޡ��쑇�N��Ѱv�Px�m����ID]���Jv��nu܆���~��l�=[��z	�p���ѣ���=�����*�n��F:�险 IS����K���"y�H�º7b=���+jL_�G��C�k�pˀ/x!5��aĠ'�D��M�eWP�*�,��̛&�%�n
Lv�P���N��ɸ��������4K3X�(S��qH�|Fe��d�fgH�++�z�w��Q1���g�$B`��J���Ur<�B����lM�7�}��k�a�MTÎ����I3�N���eJ�c��X�z�σlэN�A�l�L�6�@{z��������]�G�o��]`�]���%_>���zLeI>a��T#RN�fP
(Y|/?ie��3�AZ��Y��>��0�'=��G��s��K������S�k��hRD�7���+� ��EQ;R_x_\����^~� ��IB�) �?��?���>�яFu�9�3p�8��.���Mo��`f�q��ܿhS;-��lf�|�zb�3a� �M��i+(m4H=\<�67h����nVA���ٰ~�n��Ԍu��ӭL�x��>N��f��J����XC�h���Ry����3:]�{Yìk�<X>��OE��t�rS�a�����e8�1+H���}B~�5ہq��ڃp��q��[7�F1B�R|\6����Y\ ���y�\A��c{�SH�p+y����z�1�@[ ��N+� {p�|��d �f �2b�Bh�p�.�ռ�\��a�;bm�����\?���ؠg7��\�
k(H�ݬ���d��S���歜�����vn�f�o�7��pl�q��rC������;�c��^��UKF}T������䋷A�;�D�3�	�꣇-�R)|^���J�Y���_�L��Q;Yp��w'����+������z�������=��w�;�K_�R{���B�ey�h��So�;�D���$:jIe��{�b,@��'73��#ùS6�诺�q��қ�Rܰo����mг��:���4�`Ǐ��v�F-s��t�T �ik^�%7<�v��8�i���j�u�}�=k��W��r;`��B
�Cc>^Q>�V���E�D�*I[�
k�y���}��T�]-W�n�j����	�y]�#��V;A�6�w��."���h�"����9�o�v-�E���+�J~����?��N��R�U��ꂼ�dR
��> ��ІFhx��l�&'6�wz����-;xpq]�����'��z�S�ݍz� ���Ӧ�mo{���c���I���Z,��l�lz�Lkf�Ըa%�'��T�eyT�
C�o�u"����3�>�$jSHҲ�	�A���w�ԧ�QT:S��@���D�:I��D�Aة#�IT��J�ȳ�y6�GwIE�� �+6���?�{|������y���}�I��
����$����f�mE�h�j2�w6�9۶���0/)����I�C��½&��J2��RF9=<��
1��J�$�J��g�����S�7�'6h�i��N�Bnz�@$��V'���k���g��/<C�1ĵZU{|�U&f������z�b�F�T�6vDӱ���Cs ����f����������/^c�S�#q��-˭<#8߫E�6�^ .�֟v�̱.qW��y���'�H�Ġ��^�je��8"Kv�
�KΉ:٣O�%��Q����X}�+���s W>+K�t5R���!:#`�w��X��F/��"��8�Z�G�_.��L��#����]x��v�M/�͛C��cG�
�KF�0q�R�3�� ��<n��9o��mp�]��'.bra&�c�R�@6 x��i*��;�T�3�1�J˶l��c'��?�����+��Ѷ���`��-�N[y*����n�lO;mG\D�¬��y���ڽ���ɵM���`��d�)Xs>�]�
��L*<���'�e��e0�Y�$O�ߍZ�Ռ�xN�UNcxa�"�~��N�Z�}AVS��а'�Tt�D����1��j�XDՀ:]��#�b�0a������薆h0)q����.�Ї>sI�d<\��[����8�سx\7|�e�t��G?�����7����s�ґX#�رV>Lr�
��˃����76�c�q`d�/�`�qL �q$��mг�2Õſjd��������~�ؓ���W�������R
@�Uo��a�#7�l��������7�9d�(�>p_#�Ǒ���D�:�%%Q���8c�8�R�zݰ�Q�(>�s� �rM/�gx��:�j�Z�]�3@(ƥ� 湏�m^|Af ܇���H���dm��ݞ�:;~~������H�z��*�΀������_�r�.�|�!���@Qe^��-ڎ��؁}���){�˯��\zA��ь��F�����
g���p�
���:�Z�X*�����J��#@�C�E�|�7h�~���`�K�G��0�N��'���}�{�lv���P<���Z��zc>O�s6x��|H��k��62kw����R�]|�����-�t 1O1�Д'VH�7�+Me1�;8'M� ^Z*i�h���#hI�tC���F�ވ�����Ύ�,��*�*��C���w ��?��_(���J� �<j���/�F9v>���^�̫2�y�4�_��6w��Ϻ:؈���'��l��4��G�%y}�n:�М�!���f�9}�}�} 6}#��6�ڠg%�[J�i��k������m��>�P�yr&`C3p���pV)i���a}0�J��}��G׶V+� w�_%��^SPG���I�4��aV�I��UN���7��0�!�s���+>�Ւ����r�i��t�h-�U+U�(n��&{�UW�J��2���]�݄���p���۫���>��A ��j�](�������$�����I��]aמ��tI)j�;�o�2l�ਢ�s���K=1���sx.��=+�u���Xk.�/ʕĦ��A�<߾�бhWR� �S!X'F�Yw�+�ֲ�Z��r1�E�)g�`>�L�I0j��)Ҁ:�"��{P���8��a�9B��lujvr
�%9a.i�N��I;>�E�5��c��j����HUdP�T7L��n�q
C���|�)= �M���n�\Vy�RL�A�Ӌ����z��J���ѧ�~��]�v�o�˟^l��#sV%�`���k<&��{��MP1�|�
��J��A�l$8�t��r5����t�xo��F{��O��G��l���c�@��ԗi2���jL��QM���y�Y+W]uU/�?��)��d��mF�W1�
�� X�u�W��b`� b�}�.��Ҫ�Q�t���Z�10�1@|���X���5���)��p� 0�p��Q���������NBf�.��}�ԓRT��D�Und��>9U������9gO�UW�g'�"�[�N�����@�j���?ʋ�9~���S2δ_~����.j�LS&�����Z���m�4k�]w�]�ޫ���+��18��LF>}��k\0 
SsG�%�W�<��4�~R���p��L��t��ž��RQp-�
�J	g���>�ǹ���#��+������f1���Pi,�b���Wg ~���j��-�������㚨-H�9SUd՗�o�_��/��m"�`A����j׽�;����N�s'�����7�3 p��FE�� �H�{"��HH.6���£���T+�x��a�7虢��f��5���Vg�R�f��b���>g�ݶy�:Lj�,9)Jq�v"x+D�x}H���d� ���+12
ʐ���WN5��H��6����\e�P����7����S=MW����c�[�� (�c���L��>��z�Ii�=��tU�ŗR	3ދ��<���&�7�#�Xd7Mc1�>�&�K�i�Ҥݲ��ħ��� *��ih��{U�b�!|�ѡo�=[)�}�lwb�j@\��}��
�;1����f��)]�l�rukTE���h̋�[�ը>T)4�-~A�]T�Hă.��u,�[��:xCls�F��0;0���	�� �F�p>�y��=�*m�g�(S�F�(�OI}xG�r2����a�ޱ���y�,�U�6՘=���h�����vp�!�P�
�]�|ʞz�m���I�:c�&
�JqStPlT>e�j�A<x�	�VLH�td�6�YEi)���*�Arl��C���|���g��VZ���g�i�]w��>�b���	�\�ienm�{婴n�qz��Tд�-�I�trV��NO� f�X�A��?����TWk�[Z'��Ϝ��I��48P}�-6\��AyAh�9:��~�Q{�����.�����'�SOcF�Vc1�HFϵu�i�,%�zE={nj�Oe	��>���#�A��*����X,!�A�l���mƥ�5��۠�C�
�����}�o��O��B��n+��ö{����Q�s��:�vO.J��@q��cJR���{H���[#�9�^'�(��D�LAn�(���@�Z��G�)��8`�
����O8���1	��� mҶ�R��� ��N\��.�#���&��q"�X@[U2'>�
ߠz6SVA���$-���CZX���� [f*<�p,?\Ӓdb �Đu:�k[�ֽ�0je^�w^Z�I-*�$���b=�y�X��U��tu��OY'�5��)�2Р����uvyNЋ��|uoo������rG��V_<'����hյZ�w��B�~�Ⱦp,���#Mb�����$��?�+©�'j�zUF��;@z�6�YI��j\X�额q�Vۺ�b��ޚ�s��]v�U����p�R?�"	��Մ������5���$�� AN1j��O���H6]���Tii?a�DH��Zn~ ����V�(h�!XMt��z��v�^�<���޳c6�W_n��-�Ś�j���?|������ر� {)��HO���"�̠rV�5� ڢ����}�7h���T�%��`�mˌ����[n}~`[�a=um��67_�a�Ie&�#N��)=%�����n7�}J\�d�Mѷ����ٽ*B@*ψ�qN *�Yb�|�Ȩ5_���	���#E��:?D�{Pw��� �kt�?z ����s��f�!�e�v������	�N,�Ƈ&M���U��N�/<��\$�`%����ʡ�ngbX���Ǫ�N����x��2ܩ���U�^?��\��jh9��Y��^�u�l�F&�X�`��;��3�w�Xu#m����v�pÚ��=�$>�oV_��,P�aD�K�A��t˒֚����^Y�y5�O
�ϕ﫶g���ѫcAx���C��s�A�+���*�E]Bw�XuZ�Zu�lG9B�+� ����3�]&�U��a�p�jK�d�)�C���m�����+���w�����|�}�O�(�@���rf�����%t2B��B�op�0¦^-�:��I��l�\��˗_�o�*��Q��4��R��R�Y)h��~Jr%��,�۵!�o]�x�R�O${MT�q �g�}N����=ީ�NY���$���nB3˨ۺa�����R;���?����z�.��j۱����5�;rׯ�t��Y�~>a��A�+I���F�x_d����g�<�mO�XOb*{�D��I��ז���XPH�ة~��Y�/�?9xP�}U��X03�Ȫ�N�����rq���\�R7x_[��	臹wr��}�l�鿱���y���+���6=���漕p*��=�W)�}�y%( "@ݿݍ.p��K(�fc��}�y��(�m�O�4�7��Jm��/��;�����c~���,^��k�_c�-�1Cޤ�ڻ�~�ܯ˓�4�O},~�w�G6������W��N�ju"���G��fX�����o���g�]��b;��K��8����X��{���4�Q{b��=0|<��yU�O/�lW�>@��N�my#�h6�F��=7�XHe��j����@����6-�Vd�S�s�
x�,H���ي�-�O�V��(��|�-Λ�����|�^�����ZDZ-�]^��r5F�� ����Z������-�]�{F�|𵨓��pN��o)�Q *p%�����n���9C�4NF'��QB� ��Ԭ��KI|��+�&Jm�s��j�� ���u�sk��F�@x-�%L1=��LZ��i����'?g�~h���E��isI#\)e�M�D������ƶ��n�����o._�] -����yK6�`+�� ܩ�}l,�`)�����ʸP*���`�����a�^Oʥ��2p)�Z��T�c��I��`��*�D-�5�f��܍��\Wk-8�n���y{��OU�uߗ�|Ggx�2��D%0\ts��ߋ�e����w��'����ˌ��7�4�t�t����`��`F����n������Y#%]��t��z� ����D�2y���*�Ν�2����TT$�U+i]��˕ؿ$5K�6Ab�̅/�%����e17Mx���>�J;f���K�r�C�j�+&	ދ���jSM��_���H ��D���-u�z(��6��v��/�ZKlb�j;��bg��۪�vb�8��.8i�9cX�DuD7^�T=JK`��h�\o�r~��p%�㊟ך�{ݜcNY����a�e�Q�l��C��1�x�t	�xO7<��a :f܊�LO��rX#1�	�-*U"`x#w�_�gG���{��X�e�ڭ�u�i���b�F�Ϭ&Ղ|��LNs��KI#�r� g`!�TCT��ҝ���V���?ߊxLǈ������^W\qE�
#O��z�.D������ܞt�Өݍ�a�������'�r{r-�Y����2����Qi��C{������7��]x���X��C��7��K���:Ҥ�c&ʎ��wm� O�!��:��2����NR���.�kb�������� 5I����r��uXZ�b��ü$L�C�_��?�jfړ�FQ��=���_m��/9��^�Z�
�Нw�Ҿ��'챽Ǭޘ�fk޺j����Qc��h��<�Iֶa�z�O0XA`��H��0��
�k�'���A����7]�.�0Z���Du��k�F�J�lg�}v ��ǜ��*�' F%J��).�)L�)�C��Т�1��n��6�����x�w��gϞ���/y�/G�6�j�	��㜤� )Oe�~�m���.;�^��Kl��h�Fh��l��1=/a�|cґ�G����M���G�~Q�Nu��2����+����'+�(/n��A*3$�z�68鰓X���9ߓAx3Nt�3���#(�,
mPK,�6����a�fw����Z��d��"�i�����(id�ն=�ϱ_������7	��lۼ�fǏ�#��k+V�Xb�����P$�*�DMb��.�,F�RH��ɚ+}�c�@���7p
�����$ot��"���0�SS�5VGt:\� ��v�M7�ƞ�Gkr"(!��o*�;�������P5��ߒ�g��뮻b"旼�%��W�"ޗ�R�q��b��~�R��,�O����-��^�[��T���F�h|}9\r���,�c)Z���~�䋤c�b�l���A�������-����v*���>��������Wx]�w���뢟n�����̆y��,� i��(z_�( 0^bj�wۻ�h�O�$'��1�O�Լ��� 9���P¨T�F�w��ٳ9zE|��='���/'�ru��@Y	x�/8B�0$v��/}�KG��e[�� ����_p˔bS Z�ت��涬`��q�0����m�{�����}�=��S���J�̐��ΰ�$աc�(�Q?N:��P���J"�s�=�^���/�rs��2���>�у<!�d{����)�ͻ�~9�V��f�R�ӴV˔�?|�)+_W��Zf��"~�x<0D���6�1/E7mǪ%���K�r_�Iu~�si�K���dƻ~�`�+�8�����t`��~��n��Г$���uJ��-ñ<��#�L���g�G�17�s�OJH����~T�W9��4b��Rq�T׷�h��G��"}2��)�I�[���Cf׬�J�����w�"�|�gon$݁y���3,1l?��'��R`&Y&#��V'�jWVs���;��*a,��G����0�m'����l�D˶��;������<RD+���^�M��z�z�9\)�õ�R79��L���J]�q�6)@ə��ԗ#:�{�qn��U�P�8f՞��X�����ʓW���fl���:��`ɔ[���a{�5W�A ��x��hx��I@'}.`�\��܋_��8����IKW��?�S?��cء0 ���cy0��a�<��|�3C�/�wa�,����w�=����c&����2���aB#� ���{�>a����G~z|�R���Y��1��8�(P��n4��� �Q�
��`���{@8U��r�23���/��[� u��Ja2�ݜ�qaR3�}�n��e�}!��ϯ:�=h�ő�d����'$��t�'���Y�U	�>�po��N}���ə��ONTs	�q�����Tع$*�$jb���[:�|�[��{�id��)�r��$΅X��m}?��	�pȾ���>���h8����;ڶ�:�\{�tû/)=+ 2�06���	�.��(�mw�����k��Q5F�+��2�� 0�l���1Q���Nػ�o���3��y�e[o�˽��^���[qΈ����ΞC�Mn��WLȭ����~$}�~�;*�����q�u���9�~~:�Evm�nZ���ޭ��׉zǩ��x�7�Y��?�A/���׽n�v�����K�
?�^�8�Z`ﭷ�:탹9o`��cp>�{ؐ���
7�|s��*8�O,{�XjG���� ��r3Pzn�|�}~CJ����w\|�nL,�������7�G�%��q�q���"`�2ep���g�Y3��!�9��J��o���1	=����~f��M2WT���J��q6<p�C鯾�t���:�6v�����P��l.�n�A7�[k)[�[7QF���8�=]�p����h����r��zʠUp߭\���y�G��zg��b
S{l:�L��섃�g&���ի��,�O�1}��ۋ�@����u�r��9��m����"5�0;n�`�m��n��c���aTY�)}���D��kw�-����&[l� ����T��׋ 9�4�7��w��&���5��0 �[o��m�\��6�ݥtp�ĵ(ӃS���F7=`����ݕ�3wB���X�N�d�J��Zݏ�M�� 7`����������;�i�F�"�Hl���z9,���T.	��>���旁p �9&����Q�;�nq������4����@t�w��/D�$�(�iYII}f��er^���"]e��`~PU1���y����|B�LRC�h���kl�	'�
d�,�
0�c�-�&���Ғ;HKt����u����v������ݻ���t�=/^9�m�	g�h2]ty�����t�iAZL"o������̛�*W `��g^��l�) w7gyj�/�NR�*�<��@��P��T��!3D~�F�ϚBv`j�޺�1Q1P5P%>�&Xiky��"==VǚŊ�?��פ)2���e.�.=
gBh��X�2UҔkPڽ�NS�?�$?+�^DƵ�z�����u]Ϝ���@|� �VZ��=�I��2�k{i�����d�ʢ��]ߠEX�]#:�׌���*��\r��bV�̒`Ɵ�ɟx9X
����o�?��OA���� ��� 6�͑Z���'hͩ�3�������F{��Z�n+��S�+ƝZ��ˢ1�㼳�q���4D�q���(�VC����x�)�iB�c���(�x�����L�W\�R��ot�,���<Nn�Ml͠����F�&Mz.n��0�|v:�HJ����:�w�r1�k:"D���@7;���C���ܸ����x4q�Y6_g~e�L-:)�a�c�Y��ô�������eS��T�t��j�8�ndǇ��d�� �=��)𬨦P�h�v0��ݛ��o��t���7�������0�qݜ�6\E����X5N����6�������^mV���TL�S�M@�aX�g��J����4��4[+#��Cs)R�eb�k�ήk�B�6�� �:�u���O�{��g�p��X�Re�0F�$��5�\N6kM�r!{ՅM�?���1C�5���x�);��x;e�h�9.���bn�k��֣�!O{2r5~R��f�T�Kf�h놌�C"�����%X�i�$7�$e���&`��,��g0�^{�4u	6~C�����+L�`��` �t��m�:��al��Z�r2��Fo��G�������j5L@�$���ÃE��]�yԱ)p�=��WC�ѝO']Q�0�����`g`�"?`�f�[wh�_۠��R�/��Yh��d7�7��)��� �ڌW�U�&<aM7%(ޘl�&-���U����	�%�w��`Ǌ/f*W�'��@a@�!��+;(�
�^#cR��D`'�\���y��I�Z��ʺI~�2���r!����*���SG�y(_1��?�����o��-�T����y�SGdfХg+r�9('��9󩗳#�	sϵ,-7�l�����^�� �XTה�C��`q� l�L8_C��,�&�ՙe�u%h`e��05��Ɠ\�&����q����&���Ν�Ƭ7�wҀb�_z�F���(�!�Yk���E��/�y ��d:�S��׌�,�M߃�|/U1�ħB��^��ċ�T�Mv1���������X@@��x�K_�{���Nf�	��Wjة{��>jU�~�4 ����f]�E$\�i aDv3d&��sB�$�`�Y1/GuB7���L�z��1-�E6>�'��I��?���/��/�Q�����漊���G���ƄMjV�M��M=F�0v�YXX�L96X���&u�Ė��s�i�S���ߑ	ov�0��]��ls�曞좲�Q��zn�Rf���-:�ڰ�ONIU"���F��0j;��Rׁӯ�0iR�9�7V�:C7�R�Ә�w�^70�pV�{9��N�(;�r��4�����{���^���:�(�iH�s�� U�
�E��`�M� �|Î����V��ͅ�7i"�f4�;�j`�,�,g���,��<S��l[,-�=@��ݘ�h��g7v���|e��'��j��>&����h�NV4�ko��38�βobc.��q���zӨrF\����`ves_u����m�ct��p�MZ�K�A,?E���ϵ%4�����k���{DǍf�F���w���h��3s�����?O�*C�t< �m�N�U}+c1���fl\NS��q�{] \�#��S�z���*[Tl2r���r!Q:�dZPؚ�KD�����U���~�{�s	H��7���Ƙ%86 ���񌎘�9b�p��G;��!���3;�\-��C��iV�`V�=�W�t�y��w�!�`b��k�R���s�Ygo�EY90M�{Ӿ��^�*7�tӷ���t� �y�c.H^t��ڄ����ܕ����w�K�R�������=�
��t�y;�y{v�]����8�ԛB�`�n�)�{�����t`ߡ����vl�k��Ҏ��}�:3��B,AG��rz�����ޞ��=�q��V��9��L�^r���p&�H�)��BsF=���Vc!{�:�9;ܹc)]u�S��h��Y�ày���r����ӏn����ђz��+.K�G��j�QҘ�"�{�k�������<����5��\�']r�cz���MtG�M���O����v�����a����.��ϑ���ݬQT1���V�������}����;۷��'^�ce��j�*�ܾ3�|]�s����[��H�:5D��ID�����[�n�N�',gg�g����{����$&�:�C�ػ19ֳ}�N�\��I���1I���Xh��������+.�Z8#ӧ�a���}z]�|�h~�[�?�=��v�m�m�3vs�� ���MjB���AP�� e��Q^���s�Hm�B�򖷤?��?���w��镯|�w��H͓�Dq��(��у��o���FI��ǋa�J�[����E�xvO3��qV�j�*5�$�9��$�5���`���7�"=�9?al���*ؿ��vdlhh�뎝+&��������?�A��m ��=�)����
�L'��Pڶ��:u�E��qR�x)������ޟ����r�������}B���~K:��mv�5��^�Nfs�%����t�?H��;�o*Lc0�u������ғ�|L�/vlْZ��Y+OVӶ���߹#����?��H�{�X��_v}z�k^h�q6�:���n������O����L+X�k��	�����v�*���t�u'��c�q��*>�_|��?���j ` 5�ϯ�ӿ���O?��K��u _���<��csxם��o���j��v�];�W^����/{zZږu�uX�v�D
��߳绔�������7��Z����7���ڕk(8�� [[?���qpUv��y�_���]���²}!����o���9m`�5[��m��5���(�/~�o����-�y�^�����;�fK�s��.t���瞫R��ۇ�_���TW��yn�L�7M�ұ�l�i����d���կv'k�+�FK�L2�@9�d*Qx-B�ގmM5f�Js��������@�@ �����).�S��uf����ɍ���t���Ä�Fe�0Ĉ���E�A��ʰ��7�t�O2C:���⃉Ԑ�W,;���#�!�����[3�ܮ���{�8�y�##g(~�c� =�����Y����t衽�k����M���1�]|ۙ��:Bǘ��`�}֊��e��iea�30:�P8{q�L�V�껲��+7���g��{��ťIZƙ1�a��@���R/8xwN��Xp�_Z�Z�6>ҋ.ܕο`[Z\�}���gυi߾�n/�+�}�bڿo�m�����$j瞳�X�Yimx���L�+;L���}G�l���x����s�MȏL�䒦��/�s�X����<ώ�fﭥm��2�ٰcV�%w^��s_ ֖��=�3��ڈE�w�z:��rmt8u!�Hq�&�� �m5���`Q������Ε�K�;w���&������G�`���ׇ������w��cǢ�k*����{�=���\��=hb���d��c�K�&8V�wl%؏����w���0mhl���Ǚ��si)�d��k"��57'�Μ���2G;�1k���dSM֎"	�j���s?�s����8_�?��F)��Ϊh
%y�E|_Z��R�-X@M�2g�8��j���h���wZ>�i�Eg\�L���.��0�
fw�u�1��א��pF� ��rSq(>��F��D��]�z�� ,Db�9���w��_��4K2غ\�X�Ԑ�@b�ǉ]G�F,p^ٱ����4X\p���]{�=�ܛ���Ϧ���<|�IO~\��T�ڝBkn/���7�wpݓN0#,���T��|�[���HKۗ�EoOW^uYڱۘ�;kvHM`;]��J���T`|�onM?�����祧=�t��%�\�9Č���QV�D�����Ӿ���}S��������fl�{nK���µ~���� V���i���ih�S7|5�r��5�S��.�e�ԫ�'nӦL"���@�+t0؞�����w��}[/���������v}�=�^�Z��YY�vC��m-���;�}�>����uO�:]xɹn*@��:i?�����:;�*ZZ���7nN��v�k?qՅ�k���pSHi��2��",Uǳ���Nnڿ�7�J7~�oS׮钋/HW_uiZ��w|���&� 4�b���?���a�f�������A��>��?�t�y;�ֽ��y��Y��<T�eS��L�uwJrM'[�d�!b�)l0�}���;  �$e���ou�x�^g��������<զ�m}�(㖡��vk�I@Dx�v��=F�7�҉�[���舜*�Y2���w�c�w�d�r�25p�y�v7C�(���Ka��FdV�YV�����X�DH�Ƭ�A�N>yI���P���*��"�b�����,�}`�1�>ے�*<����=���ƺ�����ϸ:������{�Ys�0@XXr��`���rE9�y(�G>�����t�w�sU��O>+������W�pj�d�f堟��J������o�f���{[��M?0��۞^������Zc���3]J�Rv9��D�Ů}�a��?�����|��I�Ȼ�yOO��S�s�n�Kf�\�R8��������������L�?K�ݷ��ql |iz�~%��ϼ8��Y�z��׺�I�(�L�կ}#������������Q���_���o��0�N��~�f��xT6!][/��[��O�����X&�~�^�^��Wÿ �&�lnM�3�<"���q�������|6����M{|�M�}���[��7�s�s�	%;s7��ܷaZ
� t!撾��/���_ߖ�}��3YL�9'���_�~��ޅö�g�~���X�6[�ϭ�ݟ��~{�䧿��eb�����_}ëҥ�{�=��L��n�� ��l�;�\��/��j�F'?"���l�z�����Nn�U�H�����D!m�������l6�p��}9�-�Z��3p~�*�5Z>���mm�}�<L)�j�i/~�En(?� 3����R�)+�4�a\��&��ᆙA�Y��|�C4�¼�ı�I!�ɟ��������n��
2��Um ܊��9Fu�̈��m�,���ݾ���s�1��N�}������ie��tۭ&�׾��t������jKS;��Fͥ� 	�1����}���M������|���L�_��t���9�r��]��.�[�X�>��/�>�۟Ɗ�b���}0H�x��M|��Ya��	�*nO�z�uS���nL��vȄÂ-�s��>����g~#��k^a,|��q�s��hB=�ή��o�bZ��������a��ᓷ�]g>]���`.9�Ф*ܴ��Z#������_�n�X[pG�n9����䟦�_v�;��3��L@.��u�'>���?�t�@�7X�̯?~���%�=1����gɜ��s�Y93�&ﬤ[~x_z�{?����E깣���t_z��h���ڼo�=A'��,8�h�Z@��u2}�+w��i}������K�Y�??�쬍���������7��`��JkƦo��W�ܟqM-�h�?��Ϥk�{F��1O�}�͝��f���3�:�&,��)�O;A�v^�5��[���o@�=+|��/ RMt��p�?��ϟ1�g	^Q���"ܐ}YF� �F ���O�[��F���َ2L�K+���w=���ȷ���/В�M6��cp3$[���H3=I$�M06�����G?�Q�j 3�;��_�r��}=	�@�H��I�A2VU:�!��Vs�=x�����T�r�	�����z�(zg�mw����~�Ύt�}�|���~�m�o{� x�c�z`-=��aS��H/~ɥ�{\�����c܇:���0=�qW��.�A:��!b����t�}�l��I/�k���.cav��('X�]w�7 YN�\�Tcaw{����ko��>��]隧</]{��y��84��P�m���xMZ?|K"�r��NS�/J���~��������[��_���-=���٦��KLwl����-y�k��ք�!�0پ�"�d�Ԙ�iI��, �k5�}h���K��ړ�x��{�y_|�9i��a�׮����_n >rf� ߷apv�ѭl�[ץ[{w�ZX^��`���M�S�v}z��c���y�����G0ƾ�.{���os{��2]asp�	�U�OI/{�N[{�j݄����Qz�������Y��'<)=��m���*�g":���g���j,���RK���w��Ɩ�t��ķoK�{����9w̕M���m��~� |��!�2f�i�9
ႍ����'?ُ�}^����U8+�Dż���o|cZF��������	����:�`��{�= ��`m���D���iˍ3�'C���R�}�.�8�\�X�*֝7���	��H,J�1�0gl=H���8���JkH4��g�� ˎ�0�hw�)C������8�$r� �
MS�����y�����_�m�/��I�7�*o��u����)�f���$�c�Է{^Z�Ą!y�}gүy�y$l��6�!�xki۲���*=���LO���.��xW(����ܟ|I�'/4�u���.�n0�=���%D����e\�F��^}�3|V�����H{ο��m�1�����Cv���HYIW_�ܴ���;�{�%��/6�Z�ݻ.N�{�����Ҡ;p��ֆ��+�N������v��f��"c�}�����r��@���u����⍴z���򫍑ߞ��w?�g���>���i���t����=+�֧�&d�<P���g�8�oH��zz�ŏI������� ���_~��ߡtnS%�X`>���Dx哯J���-����<-\c������'�N��T^�P�8/p�l�����g��o��w.���g��;�\uͳ��������6pX.�����级>���_�YyT~k������0ը!�0�#��+��}�2(����I�H@�d��s��9��h8�L����a:w��UD��}���������@(F<�D �+;��g=��6���"8
E�5n��g�
&�����d���.��ff�X�Wǅ�������v4sB�l� ԱNv�J̋��^�Nھ��OT�"Z�ӵ�ޖ.X����O	F�I�=�H�];�2}�C�P/K�lm{eg��Q{M������3U߫XFUM���6u�0-�c4,�Jc�;���o�(������ٿ9*킁ނ�gl�ۖWҶ�(���z��⒛P�Fa�E?���"a�Z�<-~y����bJj�d�K��F���a���:��AG�3�����+9�7�ذhs3�cO�q�� �ޘ��E�@t�r���X �Ѹ�����\n;ǎS�5M��������ߎthx��υ�<#*k�vb&|�&��\^X���HR��wβ���!*�fI��{6�6�E�ڗ0u��z���p��g7��j��/,�i��0H����ǀ��	��D0c���i2J���f�q4�'�/�Kc>�7��f�JS�lDՍPsU8GЖ!��髮��q�^B@ ,�p����O|�΂�5!x����c(�3�p�IB�.�c�2�����B�I�P�Vu���#sC�����%7Ex"Bc��#
�5����F�t����sD�{, �� �08�U�v�D�t��*�]�G���މ{��ȹDכ'�g	g�VX��.j2��6q�==��3���Ң����7�j�Q�x�3�6F��p��M���9
Ï��f����
����g7L�+��լ�z�_� �v[��67y�02b>�3#�k�G�NuN
���^���4-�H*�q�l�.�q
/5J�� �g�"�n3'-P��.���Ǿi�e��+@{�5<:��ϻ?O�i4��s!�_\1�p���� >���Z��3�e9���mv���|�x�:������{L{vc��2���Mx�z^��0�%7I!	��� Б�6XH�W�=�sm�p.�^�Jj*�?���I�	oZ�[�#�b�c|��͆$ŐW�m,5b�#���/8�&�S*�G�:Ų��=G�l�_��צ�'D4Ci�¾W���FŨ;���7�JE�}��^��-��0 S���L7�B�Q��6�P&��u2g(��RL^&�'5G��r̓���[�f���L��@Ք�TA�"���ey��\^s��Y=���&��7��sX�d%Ϥ#���d�qΞ�S�F�I��$�.�!y߰�S{!�ը{���+]]��R���L���U��笻^g��j.%9H
��f�E!��Ef�9�?98�zJcAU.��Q����]6��P�zmfϹ�p��� �N��M"Y��P�&��g�7g��q�\gѴ|ϥ�X��x\n���{��)�#B�:O�����:.ܜ$�Ru<>2���g�t-)F>�0��W�x�)��r[�[zd�t�"G1�U�u!��a�؇a��F��D\�Xs<H���`�0f�UL{�uaNf+B�8畣�M�n��N�iʏ��V��*�b��t�wѝM��8�m������K�P҇$#�JI�h�9�!G�	ozϙU�+���:);_:��C���R��%|�k=�^���T��=���uP$�"��!�Cf쀵�NYR����E�i鵅�^��KF&����L�t[��s���n��5*���-s�aS��;]Pns�j���)�$|�^B�r�aO�����'XpG�g5� *z���{�lm��IE�β� � �e:����R2�:ɵu.���z.VD&X��5�&�'�v���GUj�=��hrHk	{<�Wk�i��n^�Qo�4ʢj�q!�M�CNZ��Ir%�f.��I���M��>��p����h �n�
@-׻��0�#{�.4";�N�oI	�x�D�M �֬���1q�""���QvGͽ��l�)����"H.�2�4dL�$��r@�ט�[��0!;���R�o��T����#���2���C3`i")S�i���)��M�t��u״�:����sű�5�Nw��~Y�e"�k��s<qSϠ <+�i&��穩C��y�������۰�:; �IngT�3����=���f]%r�G_c^S�x��47��*�����,CBB��r��=sM.�����(�.��Y�tfdE��6�Ԕ���$�Y�^�jf��M)�
g�.�oM� �� ��2w���E:�Ng<7��2�\���	����!�^
�!^��>�4��dVߝڀg�Xv�G6#��lLcDS�!���Mْ1+f�>1<3D�S��Ĭ������r��*�̖9{M�mU���@���p�Fs��#�jK�n�@�����~�dU����=C�EaX����j��+�h�6��eS7b�����N&7��VPPʑ�C�̒�q�4Rĕ���}�r��\X��ISƱce����*���2�z�9/�6<��Cv�?�l�g��F'��>�s
��$�G6���#�g@S!rŃS��Ռu��V^�`2]�̛�O�z'g���Q�l�.<����KN�0��"C���^��9Fn2��{^�$g��ba*�>q��J�Q�g~�n�/ZC���$W�΍�C�GwT5�N=[*����ts͸)�T:㧤e��k�*MKw֏l fDBv$��~-�[<�2��%���������C;�k�i����`g^�ٍ����p���^������n�*�#�{a�5)LD�� ��0"�̈봰H��<�=/�΂�$�aE���q�e��Ȍԝ��ȩҶ���=Kk
�tHn�$�  ��v�\wOz�o�d�����>Eo���X�d X��r���r�m�y��>F��g�ts��<8IdP���۵�^�-<��	�����٨���B���Y8"ȸ�ŉxo@��Q1�M��XgR��}�����$C���:^"?���gsI؞/{?ޤv��3|�˜�[,�B/���M" �t���\��>��T��Ft����\E��M���~t�ML���7lf�tt�y�8�7�m!u˦��x�S���\5fi.��1�{HGf4�0�]Y	�cz	��n��9���.�Hɶ��7�@PW5�u��,m����VC�y��C�4�����HGd��>��[o�^���ﲍ��,�w��^�|��hG�1P�g2^M��Fڷ�J_��_��ݹ�q��gv�u��-`�ݎW�"��`�5c���ލ�o����`��)wi��<�t[���Kw�������������/~m�T3�k=s֥��͂&r&���<c�;߾՘���!egdٰ�ƖI���r�GUӕ�������r��D�2i &g�i?t���3�MXw�q[��WK����gբ��ah܃W�릛o�݅٨��B�*W�-9h���D7�l��6ގG������ʴ����}�f/���V΀�ٴ��g�
�1�Y(r'�J� ��fW�ą%C��n$�C�	9��7�!{w򵔷�#���i����XA�N,�m$w�͔>�ZβK�o��7�?�#��B���'�Kr��S�1���Q�ěUL��l�
Q򇘵� ��$][m���ǅ���ŏ ����r�ވӀb89�=��m'X��7��8�}��Й���O��~�L�W�{熬�e�z8ruvu�PZ\�xA����� ��>�ZԒ@ƌ�{�e���}���l﷍��[nI��r[�� �9�P�N�A�����%�O}�=�>���h.�C�����Pbp����v[q�{�M\{�A���#/0��b�������?8:��uS@��e1[�5A)OB�;��d��羐r����jb2�%�=�Ո}#E��[�F�~:D��M&W�9S��Yh@���w�|��/ _�2@q}�o6{��>�;���Ye۶�Ё���jj�i�K�n��{䐔�FԬ�X����~��x4I��X�!�N�\k�Z0��=':�):b
��4j"8����S��^��ь��{1�WJ�!67Ɯ1�Gژk��K/;Xxo�D0�^�4VQ�;jZ�$w�岀S�sa�!`�c�SjL=>?���z�hS����rn��x8A�ڜ�&9�id:j%M�a�;H����ZK��VL|�uK[���?�O��G���x�[p7�GM���a�p����Mf��z����7V��q5�~{#��z��Ta��\��0�I!_ل�\���jԉ>��oz��٫aj�7n|�e��a��ٳk�Xp)��3ہ�����/ki�ӧ��X��ςU�@pv����LaD���h�Կ������Y��r���5N=�ǽp����QB�"F�Q�{��*���%�b��5?�X��GS��Gp���'�0��������S鞋w���n��l<R`���Ю�|,�,���@�Ld����n���s���]��Un�w{����Z����XSfԜ{��G��4��(����^���Rs������h�ߏ��9 �@�q* �l��XI�A3��b�0#2�v/��1d��w:!�9�ܖ�N���o���jb�Vj�!� �~�匓ж	=���ϑ�2���8���{G����1�9Nd."��w���8��j�ۼ��s,sq,�u�A�I���h�TY\�@Q8 Sf�F�L����`rصK���6��T���U\x���G�>ua�p1�!J�^�7-ƳՐ���+��x���H�=/��h�?@i3�c1�̘��N���@|+A���JA�vm5�5/a8���hю��=H���1Y9��J���#�K�e*���Y��t�h[f�֖)�ũg�ոWl�
~��s,6�;��a J�8�iB�_�x�hr�iYu��;N�p9����X�D۩�՘r��9��\�����^[�c Ȫ'#�nd�1J�CɄ�* �9r�+�͜S��G�r�a߫�x��	�ˍR�Dݔs/s<�іMц�Ր݇�(%P��TH��yl��؝�8&}��'B�[s�Bu2��p����6��.&+��-bHk�DA\����?"w��[�s�#5��L���#���b{��%_�t���qH��a7V#Ou I@��,�*�VC�+7�\}�Y"� ?��0�}���ĉ>��}��sr2��h]��:����k`���53d���8� �*��QR��:7"u�Ȉ	�Ĕ�b�\O����֖ �+=Uc�
h�#s� .%*/��R�LD^��ƹ)�@P[��XR����%k0a��8�{3q���S\��=q�m�':��$p:��cqXI;;U�hL�s��#��4 F5���0���:�I���d�M���#hSϜN:&����$�P5��Ԙ�����ܔ�Ʃ�	�`�����M��L��27(^s�5^(l�$M��q
 �&P6���ƞ
FTV�TS�8U=����z�k_�R��`��_��t����!�>��O�}�C.T��q*�t�c�j�=����od���Þ<�3?n���xQ"�e/{�W;c��Έ���/y�Ko�7g��Q  �B�/������Ee*�v�, ��(�IsO���/SEÈi�q��#�aI���^L��q�k�����E��7��b�X$�@8&PPY�E?�'=�I��Y���4I<�K�xz�=�)OI��|��ԧ���˿�I���y�s�?���(����ʝg�?��������I�u��W��������I�f����1\MQ|����E^C�أ��1������{ ��C.U�2��DK%lm�0ܡ�XJӛ��*��6��=��t�嗻$�,@�_7�D ����(ō�l���`�0�TJ����C����5,�g�a�L�����O'Oi�qB\ęqf<�" b 2&��U�J?��?�c�d ��i��	�!���gz�`uw��{���2Eo�c�; ��=�y��7���M�Ɯ�p=�6�d�N��Ki�6r�
�4h�y������IP�O~�4I#$��!�)� 3�8^��:8c'�6��1 �4}�+^�7�g~�~�M0pu�PP����A~$�93Ό3����){F��`��׿�����>;;�tXva��x!}��캊C��<���y���M|Qh���&�NEQ����sc��pq�wp�FnRࢸH
�sQ2l���xj-��M�LmF���,���V:k��1; �L2��x�~�����Z�r
%�q];3ΌG�P�����}�5�y�)Z1L�����܄�S?�S���!E:�)8��� ,��"*"Q��`�;ǀ$�XD�:��&d�����jR���b� ���L>mo��I� �0]�$�I���x!9��w�N�����i����X�Vc����[aqL.��n�gƙqf<r��%�e	^��pѾ�����zM]�g��$h��`V��g��2-D;/�rNp �[<�A$C�6���	�I]vJc����;��p�!@G�MIރ�"q���'�C *�	R�/�5;1��b���Yc�A�5����s1�?�3?�Cy@�p�p���g�?�X��1[b����L� ����ڵ�?��\	�k2=/yP��l�;�+0G�#ӄZ����t�UQ�+־�&|ʣ#�bSQ#<��[��x�ށ�2�L�)�q�|N���XP�C�d 1�)�c�m�&��_��_w�x��L�G�>��Ϲq�@��Q���V�*p�錝��83�e�h���a����T �������{y���/Т�  ���A�wԵG�l;H��bBS�#�$��WҴ����pܩ��Y�+:N߉��瞻��7����2R���
n�5���q��7ߗTSz"����;���xA�U�.�G)6�����ԣ�<?���)�i�S7�+UD0w������^o�Xo��\������vѣS�-�H}����K�������F_)X@��W���t�7LqQ�E�ٖE ��M�7'ƫ�f�2�x�F���ٻ�'��EK9�q���1�=N���M������~ћ�E��g���ȉ�Y��thW*��A�}��w)DV�7��Mnfrc�e�Ek��g�ԤF�^�;,��i���k��m~;7y̽��鎿_W['S��c>3N瘷�Ol=�e���"K�c�����.7E��oH/zы�������o�qjj�o� ���
]��H�x�j�����6��P��贿�o
�We�Z��Z.�~�u8��skn=T�Ͽ�)-W\�nP��$V�<C��&A��߀,L��~���CJx
���u�sI��3�ڞ��8��3�f#��4�̩�*��i`��������W�ES�*��)�K#�3��8]c��?�<�Io^�d��u��-N���L�����b��a�Ҷcy�؊(�=��4�A��{D"����r�m���-A�c��锹=w���`��x����=�t1\�b�f�����\��4�T�"1d�����=�d��yX8������Όy8��:����y�{�u[�W��zsQ�<�Pc� l�R4t'):�ku�83ΌS?�懶Y�h�y�8��&<�'��w�=&HH�˷���C/x���2?���W����>�'"	��>�a%��=*��\:S>�U�F�_������M)D�-���\��rp2�K5�Q�1s'���*{EG���������&�8��b�����.[N�Zʠ�j��g�
UΤe�\C��(+��f���j��jG��3�Q��B�c^g�����>�>�6T��?��� F�c�P�� :
��_��+���%��MR��b�ص�+p@X�h%��!�Z��g��oxksĠղ]��<eY�]g�L��AZ_��[5�i�t��p�ܐ��	l�HX.�p�v�vM6c�$��%6�	X�R�e� ~,C�Y��1mne2����g�6oB�wJ�0p��:�������b��c>3N߈���f�Gc�G�����T�:`�����w;�3���%4b0 ����5`�� ��Z��`�2/0�a��e9�%�q8.x�5t�3֝����~ԅ^W�l�U+sm`l0O�}uX��^��Û X_Ib�
��
�}�P$1w�,��!;���m�]~�b�T�GP-�m��)��+J�#�i#cq��"K�c����ek
�9�Òs7\�Mg��,���3��3�4��bs�&z4s��z@�}1ѱu*2WE�0;���o87��%��5@�$0�2X~���*���1Ҧ{�]������5d�I�i�\vG��	
�$1��(���?HW����(�zh�n*'^ �j����3��"@��"�H��*!S7H�5�Zbk@� l*+���/v�ü<�R%�;�1uʀ	* �1l&a�*���
o/�tS�-���t3�ٙ��1m�әqf��!�Nb�G�cq�EU^�SU>��p���'{���wyf�.˱j�@Kam�0��`�I�>Eq� ��5���\��s�po��焩�Qi	�rFk`C���|��_N?��t��d�ét��3��S 5�����_���}2e_Aa��+8�G>��h�X 7�:��ɐab��'��>�չ��&[f�t8�,�ic�PZ^��h������x#M0����,E�Y�1����pL��N�tf=��������P�6������S9A��=����L���L�G֦��0�ΜxM��暡g��Bճ[���u*���%�ߏ�i9�֔3&��S�RϺ(6T�QlI����[�T����Q���\߉eY�7y���b�����o�yf�V�<[�}F߈�I���h>�-.��0�;Q]��6�G��BW�����ǵ4o}i�D���*���x���Ҍ��Km�M���	u�͂1� �	+�-�װMS2�h�M�>���2u�NVۛd�`����>������!҉UGX7�E�bPzng���~��n<���zP*���u&���"Rڳ��c�����`�t�[V�k���0{�ũ�����d���R��U����Pw=�Mҳ���	���`9��Ua�f�<|(�y��k4W��m�3��D��6��ɟSP3��kk.cXN;����q��0DE��,"���Q��q�ц(A�s��qbcƨZ�dc�dLT�E0�wb�,�������lϟ%�d��rZ�
i����k$�g?����磹��IQ����9"��ׁ����j�;�u��p���k�5'���	J� S�G���I怈����b06���ߔH�%0)��������	�;h�C��N�8j�e�=U9�����v�^z�S�꓃���r�jE�`q21 0��=��J�j)�Z�)<�X0�I��j������l�?h$�(��I����sv�z����0���4Y7 6��v�^Y��tO�p�KȞ��~z��Ҏ�.rޘ��λ�I��E1sv(�$n�MϠ%��_�U�aH����<��z��Њ��^��o�TF[[Խ�Z�uEO��'Q�n3�M�v[=k�|E�C�MM܌�P�5��ⳬS�[���j�<T�J�V��GdB����D ��� MZQC�@=G�T��U�a�1�I�K�����c$�T�ڶ����h�k�<\l�B>J�ҵpm@59�t�|����<��`Eh@U
S�	������o��?7�#!%�*�V:�q�*j�lc�䅼h�nf�D(�ݻ�A�e)y�Z`L��j ��&H\n��b�I=5ew2e�d��L����������mS�a:�3\�����0m�Hc�i�L�o�;�L��1?$n����z]S��:�ԫ�>�*�Yl��`p=<lm渨�����.��{b~����o/J�#1a͹j��D�>��f��jck��Y�X�|Qx�"Lb�z�\" k=H��њP�n	3�(x,�{�f���	7�Pe�X�@�)Е��c��L	F��ya��9��F�>/� �}VM4|F�s]7�M;ZC�5�sH�E!x2� [�Yb�c߸H�tj��� �-�^aN�_�������7��y�w�|E�TSq��xtsD�)�d�OV��^���Ƃ*�M�t��܄<7s0^-ˈ�$Q�e0	T�GRi��q�yO���g4.�gK��b4d��c2flG6�P0 .�1f�I��ii��a|Ua��h@�En���Y/���{�nV^�s��$�z���,7f������ʓ��`>����N�P��h��L `��uIeBj��GtrD6�g��1�R#�H�&�X5jM�髽�/�f��\Q;�J�om.]s�=��hֶ�1�:�3����Q����ɼ!����(��֠��.^׫=5�v�A\x"㎎>�qt �[_�2��������K�A�F��/ӵ�=�t :�	�C#�<�u�s��^�k��jFDavl�i�>�z�2ؕȎ�v3��Q7��Ҡ���=(?�
*��D��ő��a��E�h3YZ�L���5ǖ=O\�Q��h#/��*��Be�W�lA�vX�^����~�<�*���ʩ�%��Pc-��0e�,<dc��R[���b޸g1Xݣ�����Rs��m����ܺOƑؖ����D{�
�G0��#��Jz֑-���)@����5�_	(��~�di[0�L#�D�b�1����������"���~#co3F���Z,�=�q^%����H�p$տ�^۔��q�g�&2Ui���ccp�cQ9Q�eQ��פg�\D|���N W@�-�����x��=#	�h�kk���p��V��B7,<�A����ͤ?L�����T�B):,Z���iqkB��8��c�6H���&XFcy9gj�_~�1��������
�#T��Sy���T�̀Aẜ4N��ɣ& ��Ttlsv���y�����]6�v�T/چ���0�5�V���5�,@�T��E+�)՜��(�E��&&�+۶Y4*m��Y��)���H�"�^ڂ�k�����F�?F�(
�m�՚��x���<en�YM�X�����^P	 1j�p�f���5q�<j\�b��]ku=Q(�AYj{M귀���6ؗ1��D�� k�k�ه��_p��ڋ���Ks�&��7�)��s��k���#�(��υ=*&K��f��ؽ��Ә@;lʙ�%�WLL�Ɇ���ʪ���V�d��MK����~�Y2����<�ԫ|;e��~�I �669���ML0�k�m \t��r��oRx�v~�H�$J���.a�ndw�m����[�M���juu�Ȝ��	���?7=���{|��Ճ�7�;���cr^g_��������~&��{ -�=%c2��l��;�W�������=�g"n�8X�lr���[F�%������g?�m�b�Qk��]���Cj��72�ig�V%�Mt�I�s<� q�j�6B��vZ�A�^���CmU��(��@0���2ma�� ��ԧ|>�k��>6!ҷ�76�z�����tŕO�s��.�����'n�tZ�=�|b� 	��]=��\͢\d���(������F�C��랢�"ڡ�}��s\=��@����A�	��)tO�c��?�HĮ8�G[3�aװ �ș�b6k!4�����4��u��ۖ����I������P��a�9�f���΄�Xۢȅv�����\����l��.80�;������NDWTv9��1ݾ���$8��a��G}5�cM܎'n�÷[�O�:A�c�#ۈk�i�9{Үm;�D޾���Y��i8)����7��ඥt�TK��L�F��P��?�d;��h5�}�Y�
WRJ��mz���"� O�Es�g)W}c���L/����F5��c#��~��
9��%��h�I��1�F�$��E���(� ��Ħ�&�/ ����v��J`�	׳��3�]�3'%�������{}c--��H;�9�C&K"q��c��ʆ��8d�dt�������	���}��~>Cy[�k.�i�N���=�ԥ=�~�N-�����5F�������8M5}Đh�o�i��{m�,~�mW�Y2~&���L<'2�nY�ug�Ņ�-�������w��BtDck�EWgV�����N���q��#n�u$����M�	�i�$8֘�0`g�|	'�Ԧ�T#�dݴ<�s&�D�ƺo�����IAH�r7�5�5�6�B�Ū݇��n�>V���bw�����L���Hy]���T#��V"V�!}V&(9��I�#�p���}@�]�Ҫ��F�/;v:�� SL����C�E�C�I��X}&F=�L�:Eژ��ӛ���+�w�kB���Ę2�Au�ر�E\;8F6*| <�:'v*�j���
5�l�4�ߢ���#"���8>/=1���F�����8���'q���V?z��a�K���6n�ܱ-Б-�5c�K�m����ma��1������6����պo��b�|/D���ӛ�dUiۤ�����*6�1�8���Y�x�+��U�y�LK�rw���{{Z@�3���k�bv���7ꑳ�����%cT�9�Y�Q8V�AZ��1����<�����z���.b1Z��K�f�A�ًRP����� �z:F����,#������D�Y@ -u[ -�G�G��f��0&	�s�Ĥ)�����N~��][���!�nH0a:H��0�~h��|���&�T-6�1p�%�r������N�+����T��ZN���%��69�"����qޣ3.fk�7���':�i�� �g��9r�y�}�d��|�ќ?�D�#yH%��$��g,uyq�H0�2���Tum�ox,������=.�66UՊ΂�������0S ;�vw�V�c�À�t�}nBź�)�~(���zm�~�ϧÇ�i>���n�X��?�=�DK��=����D�`����n�O���O�s�O��S�� ��qd�n�8娐�]aal6JR�C����8�8.��WLWj����qS<qt.iHȡ%{���� 5������j(�����)�#��R��_w5i@�l�W^'���L޽�,��se��;�Pdi����l�84J��ݟ�n�u���߀�Wd��J���&�����aƵ��IZ�,����lJ��M�8��h���*��ˁm��j�J�m������T�~�wƹzjL� ��v��0}�;?Hw--xDDQ�p���jºJR	�m�.���V��`ˁ1սE�ƌʅ����!��� P��Z�W�M|�}}uZ��ҶA?�����;�L�{J��ô`l��R��ᎪQZ��9�7�\YN��]��z�Kd�7��q�s���n���-A�����t���0!1FEN��V��bYb�����̥���f|�8�,%��?�߀	M_N'S�;��~�@�L���p1@���y1��1�k�u�E֗��7�2���ם���\7L�*�;4�nB{����u���0�� ����`j�"'��lmM���v7���:5����nn��A<2X���p���)2�4'��ؠ�bw�O�7��"���Nt|O�����y���cl	���W'ɀ�$UN�}�xg�{,�I����e{؛����e[#��5�T/o�i���~���mE �nM�0��RNY.l3q�ޟj`�ks6��U�R�D��y����ɚ������;��=Ʋ���� X�f�kc��&����s�6��)��Z��_�q洸�O��Y��tNZ�C�QvTm>1���L4��]�,�c!1W�d����G �8��4�}�h#Î��y�M��L�Tbև°\(%�O9O�f(?W�U	&�$0������y2���a�V�[���iLd�{���y"�a��>����l>��Qu�rB�k)fi�1r��]��m����_��1Z���d맿[�-�o�	��G��9���6o���u��9��u���Qi��6�:�%�p���X��X	��G��l�:)���56��iNm̅�aSpP��&Y�����W��:�me�iTO�O���Dc`�s&��4ZM]��^�M8��,����#���B�Ŕ�U�����h���+;R����b�	�S<����S,*߶�	�b2Cj|���"C�"@�衎!Q����~R���c�� Gl;�,#�ơ�-%X̛��� u�a���A�P≢�Wl�1m��Fk8�kꘖR�h�l�u?��Ꙫ��0���$�'o����sM�T�"�3/K�w-��&�l��Hc��N�<dGG��(���4�c�fz}�#�DƑ�b4{Ź�@|*�tsD��^0�����D�m���U<�ei���:�N7~jT��&�v�l��V�G@d�!v7���V��no�`���մ9h�#�Rj��:+���x��r�������L�u�����H�_��fd��c�w��:����9�W�"��F��v����x���!�X	,���G��s�Q��\����$�(,�������	��E#^[,����y�n�+���{�N�q���	]н0Ѧ���'@����5@�K���Ԍ�򣻝�y6��Ud'���L�4�_�I�6�T�H�GS��ޓ��dAj����Ɍy ���^Lw�Sk�E��u���(-���PG_\�c@5N�y��T�"!�^�R��{9P\27�� �%���Oa@��dRT�T��Yu�Qy|-5T����^/�ncuc����:�~ʙd�T9!y��o 	��M�J��P�G�p�I��י����kg��l;6Y�Y�hc�� 7jc6�@b��N��"��=�(���,3II�:!a�d�6L�Ʃ�6]1�*͗�S@!0�RI	�lJa�C��6#��x���ڶ�vWLmg�"/2(*�`�fo�λ.]s.�+1�NS�I6��	���2,I�1�h?h/�Fɸ���z�a53KW�
w��S ڪ��w6��Dj��Cg�$�ǹ�(N�ͯ↹�X��H ȏb��~�����v��u]J��?�*mb�*&{t��^�$p�VY�`��Z�D�����b������<1��%&��6h�+��v�?-x�*�$�� $��U�G6&�������ƍէbH���3�4?LJ,����nm��q#����z�<���
�����&B"'��D��F-7H��\e
���2[�,4����&��M�I���d�8R������h��_m�ڦ���^6,˄@�͗,�n'�D�*�=��k�����{�`�f�I����7Y�o3�x�v�!&s|G
S��<���B,�?��3d��gu�z�h#�_���:�NZ�׹w���JA@W�����>K�M�%��
LU�ak#[� .����� ��w&^d���=:n#~8FDD�SL�j�蠋�(͙b�e_>��5���I [6��p,��H�3l�d`r="s�Y*dN L�4��Q5�P� �؄��I�	��� ��-�6L:�L�w|'���7\�"N��p4L+���F���~�9'@��.ʄ�D1e�@�M�K��X4nr-T�`_�җza ���}��.�X\1uV���e��JX����[4	ިsҘt<>���Ÿ��Q�:�d
�\ �.TfpV�g�b�d4���"�o��!���Wm�x�0Pi�k�Gg��c�7�=\{z�ؘ��y�s�u���=�s/< �c����a�3�换�:HsUx	?%^H�V�39͢SL�}�*Tx��N��<����Jh��s����ў}$[�Q�E��A����V�v�C!:y�J�W(B!���Nm@a��%���4�Rf�n�*�Z)��i4��J��:9i���������q�ur4=;�A,+���B̈�&#���ﴝ[�ʄe��is��U�?�J�߰c�븬IՕQE?��MI�`*�I �P��1D��K/ubI�a�tyw��D��l�3��n�U���$g��];��Wz�>҃I��Z찡,)����{ 'L��Efx��� .��2/MX�z�!�uW�ut8Z�{Ǟ����]w���;��{�ңO�(T�~;�,�n�u�����Jc��Ļ9���F�cˈŗ2�N�5OS&��6�2��#�i�c�� <�@���vO&��?��k�d���Yp��}əyUO�j�I��[͊��ȅy��h�P���Z��<g͑���y�g�bF���h�����o����J�D/��H)�C��h���Ѱ�.l�wsrVd�J�&�nl��=ת��Z�s�x�Ɠ��̩����9/SN��Uk"th{�u`*�L�2���O�y���[a͋��U�pL̐����Dm�\1��_��w�t���������Z_҆b�r��A�=+��Z�� ^1t�h�`@͹�.�@ c�f�TS�r�0�tSD��9>�E>���M�|�3��=P_m�5Z�|I��7`̀0�O�yL1)�T�0��"���?�gΆaҔ���=��H=y��$i��E����4�>9��(��=lz�!��*wZ��o�!��p=3٢�馆9:[�x�*兺�i�ôL�1��U5%�yO宭~a�gp��r1�ln�Vؽa��k���4*5�M6�Ϯ#^��mA-nsU������_��X ������<�)Ô]8�T#@�TN�p1�-�-^S}	=�y#:��(�I��n��U$f�Ţ3�OF4U�m����ǐ�-�*�2w4n
[���A���u��l�{v$x����Mc������8�Ԧ(%R�b�k�-ΐ�F���A>��Κ���[�>'��aqi0��5�}�vHEgf4G��(��C�x�|T�b�v����e���$�b��4� �8h֊?���PR�PÆa�M�UeF�b�0:α5�t��b���Ƕ���~���'x㼃��E�쓣�ǐ4�i����dw�_��88�q��ȯMHf�O��O��O{K$���o}�mx&�caC>�M��lBm��ZJÜ=t�9��A��p}H)�4 �L���Z��rvR�+��xQϣ&(�C���c4��{�v���fZ����V�@?,�P6�ҍq���߇+[���C�l�~.�B��}u��3���������>�q��w ٰ��qb�E�K��\�8T�W�P�{bќ�؊�@o+O�l�1ck�sN��b�v14��u v�k�|���Mm �JP����t�N�mJ�FR2�χ�r��gK�� ����p�M�����][O%�b>�u_�y��.��i�y��z�F_4)�N*&����8}�C�|h��ƽ�&4X%��)�1��Nt�� b4�|��^�����p�~t\WK#=?٤�7&X0X��7qM�u�>��P��z���1Os��ԛ#tA�ⰝB͑(\<,��y�*Oi�Ǎ�k�j`�H!l��^{�Ԇ, M2��t�M�]�~x�9������l;}�:JٹAhW�υػ�4�:����g>5��{G�G�Ɣ���{�d�pZ�i���M@�Q{Y�\�,|�(h�-��>s�b`@oB��!7�`�@-�i��ձ�w��;M�[�2�����0}�4�Ʈ��Թ��&�'`�)�h�ąцmdJ�7�i�;�e�.�5=�6�!j��LE��:�1BE�]�o/�dX<�;�V�X��~���u-mm��[�&p�K폩�*D�cE�m��+�q����?��7��j���E�:��8�4�ά��-�e�6F�`~�F��ɨ㭳&�OxM�Í�!��J�]T�L}e'������\rI��)4�̚��[Qsh�6�����g�"Lt�A�mW�;���zo��]s��*�$����7�ɳQv&Z4ׇ)��DS���ֱ�U)�s�q�O%���\7?u}�R�� <��~2�Z���:�m�V�7~��n�X0�{eI��#�M�D %)�lXn
�D-X&]]
����w�ˁV=Q#x0������XY�9��`?���A�Bw2ؠz\|�%�=g�Vb`���8�(�R�6�Z�,�(|�0?�[��f���+uw��g_l����R���{�t]=����h���͹�ۻq��c9u�=?-����Ѐ����f�O�A�T6��}C��{��k!=ɀڱ֣*RZڶ-]x��q�\<5GD�AJ���j�ʆ�EK�L,p��DV�A,3o��*'�5�x���4�bW}Ւ����2���lLE���)�)�9�Z[јp:M�a^����0�8x8��ƺn�ޝvM��R�J��봲dp��!���j��!�y�!��`�~O|�h9USv�����bP�<7��s[�;}/o߾��J��P��CM �φ=�e���w<CRp���ɚ� �u�z�f�Bz<D: ���������V�4�V��4�;�U�
J�z.:c7v��b+u����\�zt���+��Jm@= �/�ls���NX�ֆgp\�6R�̓��IT,#���>,���<�y@[�^�p��|�/-m706)l��ǾKҒTɲv@��L�(;�_�C<�t[&�!5aOEV7�\%�fٔ�d3Un��̮I��,L��t�������Ҏ��Vnj ���������Â�ۢ<�p�2F�X�=����x�׆�g_�3�k�N[-�_Ӊ/�_a��h<��zի������b��y	��M����Ǝ���Ƹ���Pg-q<�1�VD��Ą�cFN�R���ņqİ�c#�����H@�{�1���Z��G>��gs}#�B�S���0��t�B����4�)��ͼ�YX`���d��VǦA��)�dߙ�����wsY�����&��h�Mh�^g*���2�u��D��J��##b4J�d���W�WݎKQ|��F�_��z/��)Z6m������1fz�&�+�w;R���=�*�T���(�6����i �Q�����������t"7�»g�]�*[1�JЈ�|���&��;y��E�Z4f����/��/��U�w��Ƅ�������Ռ��,:�x��Ԅ����,7�gΑt���"�D�v�q�^�d�n"�5^��].�=u�Q�%z�SVY�,M&j^�E� ]4@g�k��t���Rw����NZ$��>O�:�l#;����a��`�k%{��D����dV�K�7�ܤeD#�Q�����%&u;Y!F>�ϭ��ܡ�c$�W��@�k�@�=8f��d���	��O#�@��Z��f�H��/��<�ǔ�̟}so�L��\J��d�x�4�Uڜ�:�����»/ w����S�{� �N�O�7\�%��漺c	ӹ��8��8����@�<�W����^���?�A�|���p
 g)�J �u��i�J�H��	��c��M�O�9"�BMg1��`��6��K</�=n�Ȣ�jL,�E����t^}��n7��G?�̤��o�V��?�c�H&Z^q��F�͖6=���m(*�Ԩx9�l����u9�B�<C�3����^쎿�|�QAP|��i����g����,?t���qӪi�X�r��QZ�.�=,�Н��۲�86�3�̞�&4������o9K�Öp�=*\P�|�|%�E:̋z���Q���'A�.�.��-��R��[�/�4�yf�h���%tt_ڴ�L�:�K�����I�'w8I�X�g7�����L�Ns�\�C�x�.,j~ǃړ��o�Zݸ���x��,}��ż +��a�~����{i�<G�V�g�o���-F��GX���7�A�LII�-;'t�Gi�9�	kZq�ZZ,9 ��Yeɟ���1�ͅS�6Bm\&P^c��̚�����o~�g�D'���
��^���ڧ,A�h�K]z��=�n�s�$%�Λ(;U&I��p��w�kE�Ջ��zS��'^���v!��n���t�Ъ�g��Toq�$�&�y��=���-��>��1Eԓ���H���~�k���yc��s��`S���v��
��9ڀ�F�^�"�g9/�}���ϫ�ql
ӈ�&��)}?ޫ�RM;?�Fvg�����L$��g�M�lM�����{W���4(�Q�m���A�Q&lQi���%��}ዼ�e� �o�,�ʠ"����4qq��1&Ј!�Mws����C��uߟ]ߺήڻ�34���tU�}���~��o�L�͂�e���%�}w�Y�l���#�_�ş�m=?� ����;�JzH:nS^�G��f��m���꺧e��X@��>T�	��I}j=��'�i�K� F�*�[K�1.�H�"`�#�=�;-��Ս�S� �7/��J9�tL�]�=���:���j��h���§�?��W}�W����� �l���=Z�a-�*b�����P��А�I9o�sp�3$C���%v�9
6j���YHK�cx�+W�){�=��ǚw���}�io�:d��VN1a�ӈ?����5f1-J� ��u}�����8�1�ڎ\�1tP�k���ph�f���h߻`r< ����1����ZF�����@�7�ɧ���y��9�G�gl-{+4q��x�w���K�?�5l#)	��d���7�Q_����m~�����?�áF� �����-�j�Z�	�3��w�l
�E1�Fx~�NjEc*�S-�������,�������(�n�A�,�n�<�ƪC������,�^���?��r�1�1�a���@��k0�<c<�}A0�LdDk"c��D�0��5�yM�,Lt�-��|�:9��ps���
/ԍ{���%�s\ �L���߫s1�k�ZM��v�=���:4�|��=~m�	>�ȣ}Vނ��*am�o�$(����� ]��DR@ee�עд��L���M��s->��S��a�Vh߸�bΥ�+�@�i�V�㈾w��L&�X��|&�'�-:����8z�� k�ױ��(���h�=Jm�[�='������c��1]ڥ�}%������������gǏ�e���0�X�H��������{��җ�z׻�W��U��^����BQ��:��g:o���q�d$�ϩf�!��x.��|��h<����Ɂ�s� �O&7�a�j���y��"i�9}�>�:4a&:x��v�=��=%���:xC��?���q�1ji��'e<�$��j���>��p��Ӳ�r;l�9��F�h?�X�z��Ds�-?WP���1Y��QےSЄ�x�䕽�g���|ڧ/O�>;oww�L�@Ts��#uw<�Q8�_�K�z�C���!L���.��km���\�7kx$Ր���i���uԴV�D25�!�$�M(��Arۚ�j��&9�右ԧ��&��Y=����ܝ%�G�8Q4Kj��К�h�Mb	UcK���I��Ej�q���ӂ�j�7^?S���}
D� �l�%�@t�l��؏�N;���4��x��;�A��a�CA
l:�Zt 7@ȿ����1�wc���xy��έ�,+?QeNy:W�T��A����tB~��4#t��9�����P L:~��++�k�d��%l��󶯐F=��bҁl7q;�q�N��ϊ�eT��+�Ep��{�찱h{��h(�Px{�U��bqXwb~Ѓ<�=�Bq��;��Z��p�l�V��ս�����xf�+����o�����u2�E�䲬e򢂗א����w�m�L��woHmE���JE$�;񼎜5���j��<���g֒�s���¡W^��J��h�v�ԕ�;�I*�}��M�����1�<w69���4ۏ����;/}�{1�q�!�`�h/�%�W��v��3t��*<�5nҿ`�t�%T	 0A,���J��i��dMx��Tc;+� �^F�X|�+^Z �����b��H��9��z�iDB=hh�uZ�	!��M�T8a7_t���/���MozS�����z����LQ��jٞ�w^=婟��M�>O~��.���uZ�b�M�	�ޏ�&͕�I�����.�&<޽��~0j�ߠ@_�}���{�Gy��j�m8]�:���e �յ� �~}/�����ﷇ%���b*�e*m��LV�{�}�V�Ϭe�����;�ɽ�N����'}��<n������9�M�-"���֠u/4�3�o����MGM}LD�g�g���~پe�|���򓰧r���w�^	��G.<�>f��$�>j�_��=Kz/�˒����0w�F }��8yv��P�x���ȏ�HyBW��ۿ�` �,kS���Ll8�+�`]�h�j����x�Mr��K1}����i�l��F�0Ԉ��-@�p�7m>��Z��08՜h :�����9�A�\(4��_X.╯|e�v��_����Mf��|�ה8a�w�աL�t�!�Xj�P���o/IT�"�c���"���m����H����E��P���nF��{:��4�+�t��Wڍ{Q�`^���)4���1ͥ���̛e�qn��/[��2Z�N�^��j_d/~��/9m�� HH�0�8��YZ��I�i�b�2��h!3�.�k���~˷|KI�b�������_����q���Z�8H0#����#iK5^1�s��(�;ڊks'�:���S1h/<:�4��0�c6�/� �0�y_�З �f��	W���X���r�(/��hDk ���[�Z8 �6�5X�h ��6���P4�-����/�i�&&G8/N%TƗ6���(lo�y��h;�Q��+���ލY��P�	J�ٞ;�5�5����.٨�[����KS��C�:�/��m~����e;�Ns�C�oM#��VǶ��9�~��eJM�b;-@���D�Mjg���?�Lk��U����#:ɚ�ʦt�?������</Z1|1QS�IF�Xl�yL�.�n�������n�c���h���~���Hџ�n'eXSDK��~o�-��xz�9�yn����U@5�Qn�tP�����AepM�BY�$�O�tb%b�"&��m(�#@�Fռ���a֧E\�(�X�Nh�=G�$��L�}�Jj�Bo�8�+�X�o/i�MS2�F@_�z_�1&K��q��@g5,%��k��6j���tr&��[ṿ��9���~n�:�l���f���f��c���|�*R�s���T�N��:�Rt�3��"qȓ���F�3?�3P���"w�A��:d���2��5f�N��҅k��v"<ҡ�mw��s�E���������~��>�O%��s��9�QXa0G [�4n�B^����ĺA��q6�f�GkF[��a��m���Ȟ�zm���J�-��1��b����%;���(�4����h�.�6�������<���L����G�5ړ&�0Q۾OF��IC�)��t�3�U[�di� �����'�(J���SN��c\>�
Se�c3U=��{�iE��v)/���X�k��et�d�&< #��%��ǝI������'A��zqqʸ��X|뫨����v����%�΃a
�����8P��z��Zx`V!~Ҙ��h��2��f<� �f�3L��c���Vɧ���������a:��߸D?L�^�-�/��{p�H�f<�U���z�Rf���Jv�25rѧ1�b'[)������Ak�{�5C�E/�C�r���]0�H)�v Ϊ���d6��A�+�*C���=L����0�Z6Q��M��K��,������OxN�b@�H�YZ��BQ���8���F�P�_��Хh�p��x$Z�֋�#JC���fm���a��br��,$�y(��)��B�~���8��|�s�j���%����3�+�n���9�`8�㏼[֝��u��M�މ
)��P����Ė�:g}�>�3���[�Þq�E30l pI�q�ŰS�
����WO϶��%p�=]X�e���	_�����r+���Y#�qյ������I**���T��SW[q�G�s�	̂ߑ���6�Ęm~�������6܏W��CJ��35�<��qԁY`ֹ�9m`Gٔo���C�?�UN����S�=�Gn�r�͵�5�>�f���2n@$�U�m�����0����
���Y�*��*H��Kj���gL�I���Jl!�����"��+�q��Җl4����Í�q6lٛ��sQ6U,!-�i�ϕKI�a)�c�5��4SգNЧ�r���;��>{Ϻ�p��!eF=���xnk�x�*ǷU��T��y�kA����P\�7>��ris�NI�	E�@;�O���	 ��9��g֥���!:��5�����3�#�d�C�ס�}`�:�Ǉ�qR+u�T���d�)rKj�5a.@g���l��$鷋�,'ʃ�ڎx����)1F?��	���5{V"ߢY2��t�O;-{�!fK(��]a�rl��#�mn�܉�o�yE����cW�����)��sM',�4ڥr��γ�x�JTt�o�(��Ӷ=ǳH�Ů�N^��]^:��c�T��������q��,0�K�?��w̝Sr�����>I��G�N<��?h�y+��ޠ�V�w+�![�崒���~�ߗ-���4��΢m6�|: �z�W�M+<����V����!u�S�~����I
�I�$��5g�4��ٖ���rF	̫�n���~�����RGc(�FU��~��wV�
M�,@|r����b#�$ d~.�m�(���滕�|��y�vS��*�=��׶�x�ss���5�+	���^u����oAz+[yb�y��e�����d�9�xf^8#�ڱ�f�me+[�����8+�x֬R7Q/R��i7�};�3k�.�q���)�-'���<qe�OhU�^�y���*���	�N���n)H1ۛ���>{��|�Q!q�f�el^Vg2hN��5Ӕ���6_�Xd�#��B��4P���m�t[9��s|���*ӯ�`�
�O9)�,���DZ�s���\r��N�:���C$�`��kȝFΛ�h�� �i��I0�9��w�sS�3� 3��td��c�M�����='\J<��O��Mg����+[���zG1���������9��[X�
jf�X@�x�6�ŧ�\�L��CLY��j9S\�	�)'i%�����}c�yN�e�b{�k�Tw��϶V�v�=�ռ2=xUM�z�;	\3�vG#Y��y���!�o��3=9ے���Z�s/::��r����ֿ1}��`�G��Ӿ�uuz�v�;Z�԰�O�[Y�F��Ew�����+��Ȁ��C�bn��dCԓ��6<�n���f�]F_�
���� |�y�8�:���R�:�cV�����LA��%�]�o�9ۮ��vzזF��*P>�O�`O3vΫIg�Zֵ3����cb�J ���Z�f蚒L:��ӁUVU�������pV���R�٨�����bSv�����G�8_W��Q`��Ǽ8`�N�!_���`�bd�d�[�˕�MZ��t�ֳ��|�C*�������x��ǣ�2)kJ�,�L9	���]{�8�D�ʸr��IB�����.I�X��8z'���ˤiR����u�[��B��Y��ZH���w05]��������(u#����N�v
��W�."�[*3ۚ����|:m�����H���~g�8ǻe��g?��e�^��GTw&
�%.)�p��=��x�41�G�����5A�/��//�Q9�FB԰���J/�&���i��d�{M7�,̀��Ȫ���4A}N~2���� �-s�%�U�A`�
��֝+�iL�֌�ɂBtn�$����Os�ӊ��|/bXn>�q�VV������g�
l�6�#���T��d&xC�]�Q��1�����e8�vvڡ:P�}4�\L�|v���^���y����BV%�C�MHV6��8jx��g�8��]3���W}U���5��k_�ڢU��~o���		`#TB�o�x�UZh=iO#5�X�l^7�s���6Wq��-w��=��K��w�d?���bCaj�J��~�p.B�c�t�*Mv��c>�Rp�0U�jk�*��Ɗ��������+|��e��?��?-@��(s�-Q��������F��=�tI�mt� ��؎x6���lY������K��-���4��<�J���'�̆}��^_Zg���AL�p}@͘	)���v�s<��NnX����ҳR�9�4�yMM��4�$�z^:��kgIĴ�r���E0�m2��ww�I�Y�d����}�Y7�Wi�g�\��������h��'4�t�%��ri�_6��P��$:��������= �`}s}�oJ��:}Ԧi.A��Jw�	�N�CǰR����̧����R�݊���N�Gx94TL^��/yg7
u ������-��_�x�7U�9���lYM#
�4$�cʥu���x��G�e�H~�����owQ�3��e��ŹG���zCG�Pw����7�U���w����y�i�o�9_;p�x�\���_�=��X��F�<Q����;w���j�75Ԛ�Y5�7q��ǿ�����:Kd�Eܟ��`Q� N4Y6����_��%�HG����Х/y�K��P����(vL>�x�q�A��<�X�+��+E�ĺ�6�:B)��s�^��3>�h�t�������_~xٱ5#��/�Ơ4 Z1+��ԅQ���c?�cE�������5�{<q,�����tXzVW˨�ض~���ge�N6�/v�M7GlY��Lg��рp���-F]�-��>�V�)\^S�zQ6���iL���x���	��l�Xn�Yvʘ \��&`s�L�Fv�6�^�ٕ��b���^�κw=�w��)�=Yx�S��;C��E
�!���G������@�����.)8:X\��?s˘�l�c��������n�)~�J.()�$�%�[K_���
YJV%��5��?�3N_��]m�F��>�s��������׽��2�%�k�7ύs�x�[�R��s"`;%���/,�g�b ���MHݐ�cxfϷP<�>�_��]��3�\��~Y��\h/l��áŲ
 �L4M*�&C9�2��5�8��b�¯Q�cJ�-G�dr}���+t�7}�7�p�n� ��|���>�w��Ґ��W���/;-�^5;��y7��zf���x/'��k�:��4�vV��Ѽ�9[܏5�3-G�_]�X���w�����~��q�i�������4%���]:&�Bq��N��?[.<�fm�N���:ۦ��6�� yw^0i�]m������,���e���a�q������������rZ: )!��DY�?���B�o��ļ���6E����j�*HI
RF%����J:�yf3}���v'�|n2̎���:Z���Ԏ�Fay=#r�C��ъѦ�+�jX���.8N��\�F���<��4�м���备?��惥G�4�<
/�>N��4.Z1�n��G�����ſ�e C�9\�E�x��ye�i�@��݃י���ʻ;�d0�H�{������®C
p��8��i�N#�ǃ���Ԇ���>���]���+�9$â�@��]>��� �N[���f��כ��N���V�!C����u�$w8N� Iڒ����zf,��Ay5n5����C���h�Z��|9�w�n��N���]��M~ү�- @�~B����]m��=5������:��J8�981g9�t�����__@���/��|M�������=yN�%�{��9p���X&�:F3��4�
$44(N:�o�UЇ�@�pV�*؁�����}ۣ�f��~gRUx���ܣ*�s�Hh��X=��̎1\�kp]V#���X�8����1���t��_G��L�N�m��k
p�A�l� �u���ɴy���Y����On��>�\��)��J:�n4���f�j7h�,�\2ل�/FJۃ��M���#�8��a��Y�ni�䈻����W��z������>�i��d�e���Q;�l�KS���a�8q���1��d2��kq}���o~s1ɐ�]l�@r�����jS9/X��"�����T�k5U�Ѽ��C&@e�WF� �=�P���8)#��r���� ����/��������.�>	@73��*����:�ZY����H�r/>�	^l����k�q~�tD{p�i��Og�x0CC�/������;�Q��2H���n�t�����1��A�P��4���e8��t�<�q�7���{�o���sԻ��2{��g~O����o?e�\ߟ�ĕѸ{����f|�����|�k˅����\�
�:�����y8f6�μt굝	����{�m���zj��]��|b7Jz���μ���Kʹ�׉Tm�֜焳�4����O�����51�c�#�a0�%���ó�w�$}PG�lz�����ڣs�߇
�o�D5��\t�Ч(C��I"R�ab���y<������*��+^�l�5쳨ȩ4�ǻ�#r^h�!�ͻo���B�uhC���]��`ؓ������9�;�Q�K���R3���0$)�U5	����1܄I���te��il&4�<&/��{L��FE�̣%��	Z`�v���9�yN�_���=�����z3z�Ϛ��?Ҍ��E���pʝ�v����f�x������
���9��X��ۚ���m�#�q���'\9����֠8=:�|��<���7~����4���;��4�?��?o��)f%m�IY:w�(�3j:Vs#VM����F�߹�2�є�������KG��[%O$�w���]k-��P0���
���j&5���� �;ᤖ�xp14�
�bFF�E��TԸ4�O��O���~&�@�@�p���Nk�q(�߶�J���f������E;���bAx4���X�i�H]t���<��Qr�#�K�A�5	��������w���~�����?����K�S*��iY'�����9ٽ����a�했("��rOs���6�Gn�kݽ;P�>�5�����DUtϰ�<@�eA <��jċA��y	q[ x 7j������aG��l��~�fr��4�w�^�R�_���i͍eȽ�������Ȣf�+>����t�jN�vP�Ŕ�İEǄ|�� ��2՟���Q󹧑�4��,�e�8F�4�Ȑ6R���<4f�B���!�.s�����G ����/�Ғc���1>0V����x�:qG�v<�� 	��ul6b� )�����ީCv�"�l�ߘ  ~ʻ�1���^}7�19'AY`�U�@t�\��d�!�|��w,S��\jr3��t���u2��Y�o�3��/�� 1�~���^������ ݶOp��xgtown�M8*�o7�G�zFɹ�l �f;*�C���#����>�eQ����B��17�g%�n�so�'�EHl7��t��$����7�a餱�\��\fB��aB�w<�a3�ԈV�9�<��"��1�E��v7X:!���Z�GbÛ���%ݘ�ٱ.06���s�S�����^FE1f�d�b)�S
��/@C���q�w͒��J�»�1,0\K�� ~1�LfW�y��� 'k����d�3o��t��:�lR��S�0'���,1�K%�a#����?��������z����^wa�&�>�w��J�/��Bw��x�1��]�7ˊT��g���g�����w�%��j^��� ��r/�'
1�=�)�c\�3F��YF%ԭ�u�6m�{���[!�#�5^:2U9��s%�ΏԞ3�že ¶sj`ϛ2�uKԚ`>_~��+�4<FM/#C|��}k��e��mb"�����$ţ�{ؖiu�����?#e��/���:���A4M�gU�}��h����3�5h������0�B!��+�����@�ö3x�;�b��h��ۖb�c���}�� x����m��ѓ.<Dmr�8�;X��$n�JD�X�G͠�l��>��lP^NS�I׃�Q��`p_��t�f��zp��C4K ��d-�bH�P�1�GC�D[�[��-l.\-q��$`bu�
�nw1-�=��Ym��g[��ܩ@k�Q�f��iw���s��<���!�u1x��>����Ӄ��6?�aT��}n�V*����i�_��q�#�E���J�vҪ��g�#Z�z��D�tg�*��E��`	��o����A{BG��K��E*p����g|�gM8�\�
k���f��Nx�N�����r]�cn<A�;L����ދ�[̎�����w}������9 �%-�����< �/%���h��?���+_�ʢ��Rq-@��~��=Scs�_k�7=1j+�K�r���d��~���Ƕ2�Ƌ���
��
`��j��<˵����h�]sZ4�/S��� �{���(��gy�����֦2ʡ�`yέ�'����9c�gE) ԰���ӌ�Ur+�?�Ll���m>Ǚ��l2l*��N�U��E��!dFڀ�mԎ���}3]�������Ԍ2�j�M*�:8j��j��1��.)��������F�x&�{��dg������ާ�|��|�ou��e
1�B�X�,i�j~��p�,��j���� M� �C?�C%<��D
3�S���?��'&+�I.����h5��w��.�5��:Zby��?�Utџ�����= ����pˍo���FK���g�9�3�-����V���)�j�L��0I�0.+��>�����2Y�{�[f*I� �IOhp�s3��J��#�����7��lG�-?����׼�5K��Tz���$�E>���b�
m��m��K��xi�Y���+~r="��{ǳ.(tp�4���`��J�7�s�< �����JQ�?���^^Ƽr�L�/����g�'�Ά�g��w<�@�Ώ���7�����*����'xȐ�*���w��;���4���}t�'W,O�TKr܈$��YIY��~�k�,i�vI9\�p�����V�yQ�0�?�5�^ĤP$8�F�q�d��i*譺f�}�l�xUƁ�pnJXg�7&ΝP�Ƕu�:�y'	tL���	��.�i��iZ�e�#ڌE���T�Q;�ְ�KL��{<�[) ��Ǳҡ*����^F���3��+��F�ʚe��D�v�],/�;�|6o{p$	bV�B�������i�����?�3������0�LWE g'?\ +�8mM�7�́�F��1:�t��y���=�I��a�mh�ĴP��輈�y�c���%h���+�2_�K�`1���G��iz�F^*��c_��p��w=o��%�2g{�U��YD��@ƕcV�ؕ�BVQ(�~�v�"�P;M�0��a��t��r����n�\f;�FX9?�#?��Ji)��:pI2L�V	�i��*��H��b�p�n@��P���Ң�br��Rk5ᲂ�g���U��'�������_�P���P�`i9�\�T^���2��5Ip'�k1>��P{p��1=���P���0��h���6�`�4�u��VJ`t�`;4�v��zƢ��h{��}�"F٠�>zTz3���db��n�i�7�V�!�b�!�����k�.�L�̶\�ӆN���r�]@�	�x31�	Ř�B2�`���w9���y����`&�P@m �$�[�p�EN���#���a�o��9���7\.r\��W�W˸�^
T�b����厵��� l��.#��;�]�c��e��y�}�����>�++�����e/{�T*��@+f�#�5	-�jD4*�5M��#�w������YrţXƲ!���@j�\S����'��m��?��&R�?��m9���<�v(WIŴ�a�ʦ]�UTø���7:R؇�rM��x`GM���M�0T�,��5�=���Ti��J{���&0ƨ+�1� �L@��z�s�*mRJD�L��ա���=���y�UϙV���z��h�EΒ���������^�e,o0j���Z�]�\kP��0���;w}�8��Y~�t��MтKxǨo�v�.+&B!Z.��I%�C��$�����,�+\H4�����E����y�M��AZ���k��f�[��҇�;)tA���i-��I���P����n 1�;]��d�,
1Q�<�9�z�C��@It`M4J���I�i�w�.f;��Ш5a�n�!:�se\i�}e�{��P����Y�6��&xL:�,���P�K>O�}���j�h�W��ssFDʂ�c��]ES\6�՚�����3ӄ��p���3���W��ʈ��s2c�3Q��Q{GjJ���Y��*|��M����琚�����UERyO�,������W�m@�O4_�MF�a�؋�D�Mmap�Z@֬~:I�^s���r׃�����Lh<9 ���@,�cxʺ�آq.�!6���>a���b�y�ա�X��N�^�>Ԫ�k��$�/�|�ŐI7/��6r�Ӿ�p�G[�|T�cvx�2�}�G�N�p��ֆ}������ߝ&m����;A;�]���7�H��5��^�]Ԑ�� 컬Ɩ ��S��[)����T) `�A)(O���ݖ9��Ox��ؾm��Eu��;��5�ub��2���;F��
E��ǭd��4G�z4�A�6v���vz�����]c��!"�-������_������DD�������DN��vI��(���J9���c�t�[-z��i��@� �7�םE�b���,i(5d;_��E�>L��:�Nt}
P�������n�?�9}bF��`::-ƣ��8�BS�`��{��y��OV����5̪y{-�L��_�М��:7�`x��]����&�f�qK6��k9p\�LS���˘�����s�H����0�����8w�ü�>�m�'_,�Ej�#�k��r�X����/[zxe4d۝Oh_i�:6�󜩮NNk	g(�f���]���4|Q-"'�I��z���8�?]�y��U�g���}e���6��� �S>��T�ѡej4
c�N	������ͱ�bg��eb���ye=�G��e��KIj�Y��Q�����V���gu(c.5r�F|9�etD�\��2�@O�i3�ޖ���%O��h��q��C��@Q4͐�Ԇ��o4oz�p^��#��Ϛ���y�� ���i�4��K��K�c5wK��S�`�������\��2�����bD�h��|&�F�  ����ʙv�K�#�A�I5O���%��s;~�0�q
�X3ƒ�ZL����bG��[�8VoV�<��c�;q(�����G�;��lMO{�\Zne�|ѓ<מ��6"W��I�ϲ�O��
7.�b���b��ˣ�~�i��Ѱ��臅9n�,5�a�m�.� \��aw�r���e��K9��n�䖘�8w�-)��I�֤SՍi[+ֹ����\��px��"��H� �n%�'��Lx�O+[ >*�Y��{���;� �Q�[��i����� d?�ղAT�tzѧZ�n��δ[!��!7"M��,؃�1���5�1��\k$�&b>hz�=n]�M6P6��D�"�^�,<}�dE�-o�Š�6�C���D%Tl�GD�FC��v	�}a���ۅm3�I'̇�����/'��B����$B�\��E�d}zɉd�~q�p���=�p�kE^��o��>���br͛>��p���b;�|2� 6����@�����������PD��!�v�����-�(��89�R���;u �R�����ùA��C��b'�\���4�hy'{�2jkz?3�z�j�E�[T�#��Eq�M�}�F�ѣ��0���Y�}�B�y�_Fß��S�-���:= ��5`�~���.�ğ]���xt�˄:ᤗ�#��0~�>����E�r�3���$9ae�o.�KI����n`�������Ҍ���Ck9�"�5zo�Ծ �D�Q	�BU���tgֵqLn��l���b�"�f�+�#��!�����q���06�Ś$r�ir���p���^ic�ϫ�,��y���5�d�<i�����}P
�+�޴_P�r����;ݻ�'���-�佾p�Z��� 0���$�� ��|?n�3 ��T�m�v�9�>�P}gҗ�$�����C�4�A�b�E� &���N��?G����wfJ�����H���=�f�<~����3�K��>w���,��E� ��O���L:�c����\�f�p�s�#<�� ba��n7�`cD����y�~�ﵵ[w9i��]>���Z�����T�<��r|��i!��>��n�	��^�e�|���yNrKZ�A���dY��6\�Or��4f�
�6bC��i/��ݝQ��b��w�"���?���w�u����'�3k^��Oo����ь�ԁ���p�0�@������=�KʳsQ6l�qGjMFG̗��)Q�W������/��Z�?|w��������,?������I��䈗V:F3�z2�u�s§s�<��wy��Z�~!��	��K��i{��/�}�jR�s7'�׺�%�!�Y�s�c	8�6|�½���IVpN���g_�&w�?�2+��"��$%j-T�uP)i8-��VM%N�M
"���m���ȉ <ߝ��	�1�o�C�Iz_Xo��v��m�Iǭ��Q�� ��: �
#y�cް��n4��N�8�s�\{��������']m���4�Ϛ��^�	�V�\����i���v��� O�uϸ�(�1!o	��.�Z�?$34��QҔ��4�����f1n�=6o����������h~Os��f�kÇo,9��l��� �@�X��Vk	�Y$E�:'�13��u�F���@.ԙݥFc���,j�	�j�����#�}e;Y�H:0����ZD�]�<�@&���t��/J�┅Z�BI�vͬ��\H|9Fe�s�1}&u�d�Ny��o���8!`6#'w4�!�)�|n��q������C0o4و	���`^���5���;�+��i�;�=�u <jw�G��7����o����G3��x�B�̺�8�+�;�3��<�#��֯Q�yo�1�='<ҟKi��W���qs}�j���,?�9���^�����Y?!M��:����	~5P����?3lP�H�tq�>Qs��djvu��<��J�El�s'H:�k�C���j�ׅlՂ��B���Ͽl˚]v�Q�~�����ĢTH�����\��K��9?Wj�w�B��4rr)˝���˻��VM�H��M �)���~q��d2e������}�}����
�ģ^����op��Bmt`�N̄�=>lf�Ǔ��mv�����G�R+�x1���f���
��;K�[,�s�{�f�=;��w�i����'�&��u��i�Bi��Y������8ps��䲉�����f� ��[J��Y���L�o|�hC��vI߇��{�+MZ�	5/�B�8 "��\�l�Զ��_��"Y�~��h��
㣎�Jg3�vG��K��M��']QYb��E�1�]�m�сK�7����M�aP���o����(�8�(��!	��,6y�^�]��i�;AH�k#S����D5L�;E��ܝ�N�j~v�Z�쀁Jڤ��N��G�C��I�7��l�[hD���yoëa^�O�JUƄ���3�#�ݻ�v�ּ[�g���M:�e��B�Lk0犝INZE
iS�\���F�Ms�|�n��H�I�$i 5�z�y-a?�HB��%��\���+;�����.�%�8�|������9fy��M�q�9�.�i���RY�]��x_����N�����H*��?Z�Z�\�S��R舝����qK��x�����g>�����MG� ��>��>�������	���Ex�z��M��'�w�]5����گ����4�ɚp�{s;'S��` D�:��o�S���v]с!pg�u�2��R�� x��h�B;�Hs���=�Kl_�lT���;*�w���I�N�E����vJ!z��I� s2���}վV��&�hN��$Qp��U�e���,���_u����[m�;��&X�;��L3������,�z7��zK:�8���g�{g�*��R�|�צ���5��`{�Qv����tW�a��S`?���
ճ�/���M�E{r 2�a}��=�䗣�R��偭t�dc0�͢!�E5/F�d@���|��k�v�-��}ٗ5�����R��S>�S������y�4���I�pߑ�i��'�)`6kv�t����$:���������6����N3ݙ���ʼb�K�q�媜7m{_簟sS�B�m�
�/F%�uP�.��,�:��R�S���2���a����i5��&D��I-+��UϷ�=]Xұ�.���;%A�62�$�$���~�Gf昚r}Q�I��#>na8�����pQ�8����He����X��۫�i����2�aB�)�d�L�y>nK����fo:��N;\4����m^���u ���D@��Q��t�uP�	UbB+6p�m�8��������������rr��. �M�m���B�,��Yq��Wq���i�;m�A7�4�����.���%��D�ᜦ�{�-���=M�h�(�[�7���^���34��B�L���g���M�U��i��U��8`O0������o}�Ȫw�%��:�v��V����,���*Kc���m׋��'}?��Ԁ��s�����)��җ����H��,T�wql��
�DBsF�d�$wJ�e��%DGt��|>k�by���^3� Z(+����̔!�A�3�*������AU��N��1Qu��hK/1�x��P���_~SQo���Tۏ��ਜ�j����̫�O�����Ng�����o~�E{���[��:��;P������������%�4U�<`	8���;8������B�4I*ƶ'u�Be����hĀ1��IB�B	g]xNք��j��3�ǣ^�EM�Q��}������=
Ʈ0�4B��3xd�EB�&�AS)�J�~��_] �M���Ƨ1�\f�1u���[��ǻH=AIRnոv�/���7��^���BD��C��98� p��Z�d�ִ�����hJ?�B*��	㬫�
�ˠ#��a��rŸq�F���o��  �8IDAT<�Tf"ځm���0��[���#�#<�+�u�t�����7���s@@������r�g}�g-CI|�4�.#Tf+[�ʭ*��|�(k�����1��~�`8b(���~"�=h8l`�N��p��ɗ�;:s,������I�LZ���7t2j�%=�{�:x �z�]@j;s��Y��Pb��N6VW>��>8����#/~�~��m8�ʩI������l�NK ��(���r��}�k�e���5�w�,�T�����"�YsM}N��3�;P�4_��k ��U�$�����9��\x�p;u�(���7��~�}�'�:�������Yіm(x^�u�4@�W Z�i^�"����%������s�G�u��	��2ƶ������܇�D��bf�z6 _АZ��V
x�N˄��`����%�ŀ�5˥22�c�j ���,
���K��&��ɧ���-/��ݴ�_�E��G�kK\kF+���Z'"y�	�ѐ��Фx��^V��[���Y�X�X����7��7�r��l��9�7���w|�w���/� �@x���%��_���Zǉ-�&�
�%X�ߌ��c��L�87&6�
�������	��S�_�҈W:�,9�ڝ\)���X����I�z�Ь.�+�aŒ�5��h	V+ N��<��f��ߒ�6���[��V�N1�
�{��{
�����/�b�-�jf�~z�DVN3٪�H�6g,�a��>�]{-��gC^f<N�����S��;���N�"܃���馂�1�j�� �4�2�����_����T���%���|��}]��w��$f�[Cs��L-�bH���L��<uH���V�陕����.q�Dc����J��������YW[�P�Lٖ"UcN�0����:8Y�,���>���1[�m'��A�ӄg��br6k��%���],_\�4r��Y�%�=�43���2���46ǲ*q/�l�]����5��R�[�V/�R��W������r�ŰS��o��o]�����I?��?\xa�1�ŐUƳU�bUVf��U0ӿ�gfg���h|�i���|ҩ���4�~�o6_`��?�c�E����T_�H�p��2كP�Cd5����IK�	w�&�U�LIEn��[H���*c*�"wB�me+`���"�o��-�up�8 ��1�82��v-A,q��\�Y�ĲL'g�s��6��������.�H?��фǋ�f��7tܙF�~bfn��d����0�Y��!���;���<�aú�}jv���G�c�
	�:u�2����h8Hub�m�D)����W =�������:�M���`��q ̼c��=��J��
^bG�p�ω�H���ѩ�d>8(qo�A�b�2�#�������.'1 JL���^J_*�T$�1/ $�wӎ�C�')�/zыJb�;�����A��?��%�.k#wJ�F�$y�e��4���
���uի�l�N7�k���ې2/�~��?�ap�}�H9F�Cy��%b�,�Ԁ�^�{qOl��<�E�҇T���9u� <�L
'Oˍy����J�i���������v��� ��FLа� jf�$8Ǒ����庿�+�R���ჸ�O��O���[��vq�����z#�=k�[�\�$%�8��.h�#j�y�o�v�c,`,���H����g^���{�W��������*��C�y��=x�&�3�����Ek£�ɂ�����;�� �GԼ�%/*�����Z�&i$�<��/G�9߬:���9נ���C?�C�Ꮉ> N�Q�Z:��ِ�ŝ!��N���mk.[꺳��1�u���lǭl�v�������5b�`�%m֬�e����峟���(ו�����k<C���!^��6��]<'\d�� z��~�l"�����R��*`4/'��Cb����2��|�;���w��h�hŖ�C�u���3�3���@�u>5��'��� �I��饈N���[�����ϭl�v
 ����D�*�H��IOHk䄶RR�ϠM��Jk4i	�Ȑ�/�!1��#ΝA�l�g�XM�ݖ*���}6� �����/��n�����aš6DF �2 �/�JĊB���x�;�F��I 2��r��gl��w�hq�9Y�5;~�6�񻹘}������s2�7-,���=ϩ��u0V�#�Fw�c�N�,c{�ql�VF�tv��oDQ��qj��o��ͺ�j�uq���V�������}��ssN��E���ķĮ`=
%�ό��1���=
#�FFP�E�"�5�%����e�V6iܿ޼�mo���tB8xV@چ�Ù�j��􆚜D�(������K��`K� br���D��u2����;�7�r��sq�kC���1�.|Zr��c�tp��ǖW>Y쟌2��>5�&��C#mr�U���fƙ�Mnt���Y�ܸ-ʼg�Iw�B-�*�?�����'�z-[���8 L�b�S#���kv�\������:�g�t�u����l����?��#�[���t�E�<^���v�蒇DtX��J��a�!�u�B�X~�Ŀ�:Y��8x�>G�mp���p�R&T`�3:�B��Ӟ����;�io��a���0���$˰
~��c�mM���m�̳�U�;�ᣵ��sX2���(�˦��+RR� 1�Nm��;� ����	��o\Ì��C8���N[@JCw�`6�u6-q�t��6�z]V���	��4_�� R�_~ZH�0���LM
����?��>�Bl(���S ����Ǧ��h���)a���$˪P�	�����:���83N���[��2�O���'_oi��ՒTD����C@�Vn�ASŇ��"���.�ck�Uy��L���n�P�V�����P*�����r���v�1�Yˡ���>�3�Մg�Cs�lO9��sf�������QhN��fϹ���P�P�"�/���Pǝ+:���,j��+�A2�G�2���Ƴ��L��(GԂ�ГRpR&H��jBjdy"OK��vK u�d��mm�Q����8�9�F�d��}�{�of���;��P����Q��,J��q���2����
��#k�Ǔnb�݇�Eg֌8�8�bjV�F�\�n���P	��Eٱ�������F�3w;�l�����d��YR�uPІ,2~����`�@����ȅ���\͊���̫�3��]��'����r�d;ٞ��Z�i�G��s"��a
 �Fm�
�^W�Ns.y�[�;��U���cbP��!���$~^Y�&�|s0T�o���&�/sV�ɲ�R3e9)�Ԩ����N�8�&#�	W�1�.��!��%s�����9x�^�PVQjA�'��馆�3�6k���\�j��EZɶ�|���C���%WK�'��ɬr���K��y�_���r���s|5�#�A)�2!���5	�i�;U����4��R�]�R����Vd�^����m��~��_��(��v�9��`������t*�J(Hy��k�����t�X�����8����U�:	�j�`�8��LS|&)��RMi����F@\)J�E_�E��=���_�Ņ�$�	���>j����ٟ-��'8�������O~�G�p�ܓh�/��/)�d�
R��>[�q<B��ù8���?�G��	M�Yu7�--s������\o��*�-����F�i�;����9��V>Xƨ�C.��'�*0�O.�����$~w^Y��o��4�\��t.�1��̂�h8��p�2����㽒FpM*'c/�(\\��<v���J�p\^���w�� +٠�����Xw�=I��ⳟ\��c�[�1�a����'~∖Hb�ԡ�������<�9��#��ׯ��M�茉��a;��՟g[{~M�&�+fy��A�\��+�ͳr�浪�k9)S���M����k��e˺{��K>0=��<���Ϡp&h�
��L���J�w�Iih=x�4�r˗�����i��} w��2�vff8���q��X0�S��Z�E��aI��ß�q±V1D��c䀴�kh���1�9|�3�9�IH�c�A�A8�>�$�#���	�F�
��!}*z:Jk�RNP�.O�D��l����7�Vk����.����t���'�"��QF� �9R[�~�����{r.&*�I~�~C��ⰽ1w�(ը�q���f1~<K�;mHf�UZA�*�Nz,��m����IL6��	{-�<B]�P}����w�w����k���; �FIIYƃ�gL*ڷ�]2��O��1α�c��ˤ���w����H^���s��+�z-k��p
I-�ּ�9��Ԁ{���y:EM(� �4��Pe�0ǺK,@�Y�ɑ< }ҳ:�QKKm<�ޘ������[�*9λ%��2%Cǵڙf~�������~D� ���G �L�1��G]&�p.�e��yܗ�\Is�9:c�ύ�ВJ�t�j�Y���3lS۳NF��͘�\(<&�U~�S>��o�����Z�����*� K�S����.��v$�Y��EI�Ey������('�geC��s�F�A��	S��4M����-	&���~�`�4�k��s�A���:�z�5�Z�C2��.p�v+o�5��0����ukǩ�K:˱!�����*�z?�,A�E��������V���Nj��LJ���'>m�u/:E�b�7��k�YtrH��>Y6z�2v@���1�N��N��V�:�x���H���Ni =�H��1	�|D+v��jY���I���#��W�hz� �O�x���x����xԴ��2�;O�Im��ԨS�κ"��L�3z^��˒��6+7_W�������]��T�VaIM���*'^Ƹ��k _��%.x���Ό�'�Ho��7������\�O�o���E&c�0�:���8��PA��M�8���G\�8�D��ƩV0��� �1�P���t�5��L���>w,q�z-��'��I��*�OC`�����9�)x^���B�b�j�� �v�SJ �tw�����HW�{�3��g���4�l:�\rK3۹�z��<�ݥ\�l����E����OG�ٸnM��>H�8���`�[x��ɚ�hi��t�|���ef��	�p���s��UrA��v�Zc�T����F�{���fD%q�$@L;F��3� �"'5�V�-����w���^ku��U+���T�L�������2P�E��L�zQ�컼�3�OGlƆƘN�|���ZWY^���w�s���B. 0sE�2��2��4~��Oȅ�~�����N��'�����4���v��ݹ���{��r�nI[p	"�2/d�<WhӌyA��QIM�I�LS����� Nэ/��//�������'b�d]��$�Ok�KG+���ns��}?�>ۛ6��t��-��9�)��Pg��� ��D�	��������` R�/�K�3XX�X�l3\K]��JC$հ�$�w%��ꐷ\ 385�4��G ^e�
����ч����>�<A���@j DRK��p����XJG~Xm��E:-)�ia��-L���_�y$�`������K<<�s�g|�{�S
�[�tM�B��^Q"�S?�So��N_��'`��F��]�\�cn�mG�Ō����W��> 7[6�������/~IE���ښ� ��S����~����J�4 ���w$L)����%��/���{��	�����e�y�M7��r~�Yo�B�/9Ư=�ؒ�-Z�@8If�ġ-�R�Z����'�������>�nU:��j-hS����[/�d�ߵT�.Gj��P"�Y���5��x�L�I*$��y���~~������!iiy���Tº9ʱ�!衇J��ׯ}�k��ء�q
�K�x����QI�^�E|��F�7(@`���������e
A���x9 ���Z�A��r�8�[z�\}����>�SK�#;k��`�g����|тY�ȼa%�;���=/%��r?�Nxӛ�TJ(�n�V'�|_�_P��k
�9��l�U��xܛ�A}Q:ig��r�פ�>��?=R�����se�E�J$��=�yw_ϡk��ng�^fA8��4VDS�v�n���gc@q-��o��� X�TIJ����N�MP^j�`���v|$�'�@�@=��Z�H�@
C�Pm��pN�ǉ�%&A��oy�[�_��_+������%��X+0�(o� ,�E$�0Wğ���^���<P��^h�(��/��pٸ���&P)�1�+l;��M�Ox�S� n�$�x����Լ4{=�>�`���K�����<���/��/��|ei|�C�(���ȁ�N,�!��9�~k;^�nǤCE�L���8�a�����2#�`zd��r� �9��^k�h����\׺��,@[�<��Lzhk7H90��Eӂ3�,=�5�Z��:�2�;�65b?CR�^E{(*�akc�:��������ƨפ}��Ѐ�!N�3�s��{���s?�s��@��uH�� �@�{�mso����ŌfЄ/>:b>oG�Q;�ﴺa�y��>��E����������ұc\�������.Z-ׁw��0s`���W�������������u�5��ۿ��vr=���`�I��1�-�Ef1_,�Y����>��`���W�H��m�sZ¸]ہ����:h�<��a]�WϺ}ķW���x�+
 1���hY*lO��0��p��HWq�5@��K���\����1T/��T��	|x��_]ޑ9��7�qI�!���! �Ջe���i_��_ۼ��/l~��~�Ȃ��8ݠ `����Y U�2$�y(����;�8R�����^�L�I��:��p��Bf�<�'�q����bGs�Q-�FD�G��]�h(�;����
Au�4�4)���q�#��'I�tZ^���[�����ɖ�v��mM��l�hLLV)��t\�Wڅ�-��q�il�[/9�����4]M7	��0�|q�*][��W���	���F�6���^#�?3��Hϫ�jA�q���ь��]7G9������?+`
}/�jz�g�*v�Y�g��B�s��SN���P�xVh���������£#J�·jF�U���"X��qGd ӎ����P�<y9h	���
�'Z N3~%�/��\n��},��8�J���&��`�rq��g�.u0�q�d�����m�3=�I2�����dMm���{�+�fT���ٛ8'�r1��9�%��@���1� J�/�̾7�\^�qa8b��9�~g�U.� �1�>�4���u�k���ƍ�"�	��������jhj��,U�r��bA �Rp��4��d�{�myN~�b�9y/���vHŅ�΀W��^�aT��Թ���xM����vԍ�7�O���%R�/��/����� �أ!;8r[mX�I�ՄՍ�	��c�p��ꒋ1"������t�����!W��˭M��צ]���`�M��}��L+A 6D-���5���9�����x߭�:���e"��$����XT�
C>��`� � ���k��q�5���Z�
�s�I4�S��sƏ�w��~'���m�F�M�彩m̽P��`�u���=$yӥ}�
��O@5�����5�p�C:�td���� ��f�Z9D�ݳ\�&܎ǋŌ������%yHwS��r���ꏨ�f�$�J&�/�@W��x���vN;�ḁϲI���X��$�L��<Y���Y,��4j\�;��_?��hP���$t~~��T�`5�w�����$Ƿ��/����C��U\k��wU0��r��ߌy�_p�������,�c|y�t�^ř �o�����Q�Q$�)���D'�ǻ�.���,�/?mCA�6b�ءu�����}M���IR�`,%��Y+�Q��X0b��3�ɚ𸃠Yߐ��t��/6��4�SK�������CK`��R�v��0� ?9^���gpX�����zQ�Y�<��\�.,.����`)�.L(�52`~+�#u��N4�c�Ɋ���N��ܼ��� �J�;d�QFZ�^��#�d��?F�V�L�b�G 7�%�@��e�C�N�x�Q8(@��M�1�y3yV ؈��`��}w?��:-���W9@ՄYDT�2cϮ��Ԁs2Oǅm.qjM�ǒ�WV��<���e��ڹw��X� �+�����?���\��\���fŦ�����^aޖ`������,׋��]����}D:M�m�6t��5li'ʖ���6ʶC(/(
�UyWw#G��DH����43J&3��Y.|�Id4����^�4�|R�D�Pj��9��h���-�R���f�$�2��:�8(�����k��۾� ��~�����A��$�+��
O:@]��R��`�-�
�]��7:||<�`O��0�:h`�Q��R�e���f���������+��e_�A���(��� `��P3�s>˼yM�;Y䆙���&j�f��r�:<՘�����r+�+iN�4?1�	äo��˘Գ�Z�*mڟ'��B�T��7p?(�l	��?s���� -�3︟<�ڦ�8�7b��!��I�x��Fn�u��E%CF�K^����n��2��cwIg�JMǩH&Xg�"�[Z(����h���2�#�N؆��E01>����_:\4R��d;��A`�[�<�,�#�*�*�i�I=����Ⱥ�C4��PB�<����|6_:�)�����M�IN���{k	l���Em���(c葤ҩ�<I�J�	�1;�8s���"B>ǌ�F�.U�5��\���u��h�@F:��D����9o{��ʻ���>����P2���]��<3eP�W�+��j�$�����g�3��L:�J�?��c�D>���IZp�fzVYi�?�>�-�
���IEh��j�?�L~�!<0Vd��42���nI@�M�G�Nq�����=�@�=C��`�� �3������6�e�7z+�#�8a<耡cے�I���* ��;rHUf(�	[����w3+O��s&���q�Xs���*�������KA�����N\'�$܋g{��87���L�������,�����b�3D��YT�Ѩw��j�b6g�l'��h<-�0�>*3��?��J�����Y� )�j����rMz=��㚬pi�	@\�e/{Y�Q�F��Ȭ�Հ3f�,�W���������P��uO8���(��*���'��i�M[�3DK&)�4<J8�ag�(>g��%�̶�?����1����jق0���6��|��*@�ʔJV��Y;ƨ�\�|דD����zы^TƸad +��Q7Դ��-Fy�y~�s2輇�6-m��E�� '!�p�>r����k�	�%��N��� �>�����q�16.�A�`ry)_F�$7����А�wr�v*�!�y�k��C�;���0��?�S?�ܜ03��(M��e�y��̠2�Î7
BK��� 1aP�`�Y�t[�\Y�	�L^�P1��΅$-!�M�C[�\��Q�I��r[$5W~瘴l��� 67x徆�ɍf0�OJ�N�� ~9eD�.��8� �o��on|��bU�) 	�5�_���F� ^p<ֳ�������Z���%X��y�p�����͞A6J[��R:����L2L�O��Oj^��7ׯ�h>��?[�4���1�P**�����dU�=�Ƥb�����\)%G�Y��%7�xa;T�G�k3���@����9"�nQ��J��7*e�W�ˊ��N�\�5!�Y�G�8,`�NS��K���[���%#�$�o�"B,�W �����sė.�A�2 :��GY�s��	#�1p�`1GTPL쑣U[�Ӥ�zj��=�q���|S���Y  MFYB����u���
j�0������%>ڭ��ƿ뻾���;���e��1�F��rQ����,���r����Fb����5
^i�̦VM\����LZ�����a���d�����B�JY��O�����q`����6��%f���T&~�`��>v�&�⬐�X.iBls�r�i@;�lp}�\[���5��jIj5���8�@|���[��!���B��5r����A�t^�Y.�~�w�c�t�E"ǔ\*���sF$�J{dd��ajZ�|f�7c׹�U�)I�<+`��=�,
�S�V����=`���������u�ٗ���<�=�G#ϑ{?*�M�j��0�'�xtu�����_X^�	~%�Z ���Fc�Γ��@ ��uY�seup
�TMm��1���s@� �^�Z��Y������iz���j�i�aj���).Vj�75b@�j_��4uP'sMMX�~�1�Y_�- ���7���R���&�dn� ��s,�;[j�9�� H�$����AQ@Q�XY2V�_��Hh	C89��uZMe�IV#�|� �r�(��םj�<�s-B]��rĵr6�0���q����9��a�R���RM/�h~���<�h������bL��#Y�So,�Aʳf���������4�\Y�h��O��2����߮�6��(i�;Y��u�����Tn�%��EMg����E��4߭6|�Z`~F)V�m�X�:��R3<����  cq��q�?"˛r� z.�)�����e>����DI�5����\��ID%'��8�����7,'�����gý��wJ��1*-Fx���蘗�U�ח��y�CX��[k%�yoF3t�	�3q%�B��.��8�Y����W�Q_��o}�[�g�z�;%�Y�p��Sǂ�W��;��;CE\��m�d�K�!�J}7�h����!���?�>�1Ъ���-�!x� ߂��K�iMI�S��T�b_e���r,> �հDnnmeqr^�%�|�'�����ź��^�X3�6钌D�8Dʄ��[�%�㴐O9k�q,�<���:�sg񌭷x�A�0Ϩ�F`@�oJO��j����L�B*�=������7��1x;Tt��̧C
s�!ӱ�(A�����6��3�:�ģQ�D�z1��a���d�Ϡ�SNX��n ��q�vЛ�o8��9�,p#�ʨ���q�p�[	w���Ο�{ Tm13��.J-1N�qo|-�`h-�1�8�9f� (f���%c-w~q����_����n��c�z�'	mF���_���/��k[a��q���A8,�:X�?�EF����+�˱�k�$�������x|I!j8�\yv&}��^�sZ��+�������%����-���m9a���@q�M' �j�)ʧ���}�<8�L���Pc�����Lj5�h�	C?p�Zj�m+�c	��Nt���'����ݿ+��$p��4�jpy�:
�I�ǹ"`"����%�u9�,6��kX�Q�Z�>���~��o��r]�b���vQYWV�(Ƴ���F2�X ����S9�����` �)��iY�FP\��Yݝ�c���ɝfہ�������`r,A@U^�%M$�a!�& vb��� ���}�W�t��ۮ��b'Y@�Z�f5�����t&X��N�೚�C��{9RO��Y0�w�&
?L*�+�i�,��:�>S�SMm/�8X:�̮�Tz ��,c�}7��3��g��vN�$�/Ǡ�RF�9XN闬֦��u,�mq�,��s/J�I�A*ù�iھc.��8�xN��N��y� �Ĺ.��nz��>IRz9��,a�������&�ф�����軓%#4L�*9?8q&�+sZ��[�X3��)�#ﵕ��U���p�Ϛ��@k�&�"�R���C�{�/%?�|5O�RƔuX�_��{�Np�P�E�c�C�;D�X�`O��Ys�1��o�[`F?����*`f�|i��'��nV����\VY'��(�ssQƣҿ�ч�H���uWb�b�fQ��j��R#1[��;�ZD������V.Oj�A����c�!�t@��zr��
��HM1��R4�����ȥ��G����s�i��ؤ�q�=�������1ƽ���:M8ۢ�<\���(�~�����*�Z��(e��C��ƹ�dg��]܆9�(N&$'nz�kn�E*M�Ui+�:�A�OXT-5��H�B�֨\p9�T����:,��@̤���\�	��Ka��
�z�9�D6�Y�T�ۈ	�I� ZgY;Bz�{?���=�(-��Ƽ��P����2��q�^����c�&�n��� ��C~M�;�6�E�9�
�#F�j@��A=8�<�֞��VҏwI���-��c�41iUHZ�u�0 9F�u,���Z�TcG�㽾��ݑ[N@�FEj�n��C�{fVYf�%���]8�gH��\f�'�h�7���n.�g�� ������p �5���w; #�N�Bm�d�4�2?�ZH=�:u+�'�8F�'1�>�`� ������4r�[6��u#�w��Aҁ��?������+_j"�[()?ñ�ְP�Mm^P`��z�e(NIH���+�
�Wq��%�h�+5�Kq̝Vj �H�U���� ��Ť�T3�����ñ`VyJsP�N���H�' KG���/^�n����yV�c� sg�?�O���cܬ�5��rH��2�<���&/�q(S��2ؑ?MFk��*,�`|�r"/f�3��EM��#��}�� �`��"߭�b�tC��sn����\�V.WrqK>���2��H�7����ke�ǆ�R֞6�غ���9��v�����@VU�y�ȵ������PM'��s�C�;<6kN��:���JXu�Eʺ{]�p2O��-屲�1w)�d]U3�6	q��r<mb&��5�g�{��I�d�a2�I�)�U�����L��&��ˑ$
?#q���n�Ԥj�Q�5ـ1a�+=���6���ƕ#��qh��,Uh�E�.˙����sezr��Ҏ�t̩A�I���6$�$	������Eh_\4W|�ս
����6�4�ɸ%A�d������ Ð%wp���.��z@Mذd��9 WZ��U$�]}X/}�KK}
��	��Q�p��ʽ�61UD�\���ǥ*0m>��NI��o���/��|�V�c�=L�ɰC��^S.?7�o&��l�1`�	7�x����W�$������L4��*O|����
�l�U�;�l�[��)�Ǜ�f+گގ�	1?2Hm��'Z����~�k���e�;�ȝ5���*�H֡ �~��8���F�P��1@d�7��:/���;e >��3�[R���D��hՀ�:��G>�4qd�L�����_��R���g����4,/kf : 3�ٍM]��/]h<��f�fX 2��u�S+'���h����P���O*{��5ݐ�+]��s�� �i$�kG�O.� 3���Ea���u�+;�ґ=d�x�[����/�r���^��ׅ�$Ȩ]��ec��z�q�wX��k��֯�t���B�!�@�?���`��SǍ��u�Xx��q9���t�w$����K�dD��R�H�wr�逳�+0�u��3N��05A�k�E���o*9�Z�!o\�qc��J�*m�~G��̴h��X���:�d|��D]bv�aAr/F�CF����h�:2"(�Z����Va��#(4�3�E���g6�IJ�~PЄ��O�ce-'|p���C��bC��i�Xn<�	���E�ç��{�!��f��"/(�MU#4ƕdg�׽���m���7ӎ�B����z�j�j_f��~x�x�+W�݌;���f��3lĸj+��+y�ޔmۣ!Grq��j<��I�k���A.F\ۺ���1���ܚP.Y�$(�=���M�w�x,��ϡ{T�=��I;��G�8�������~��e����sj��t3O~������Sk6�LcK�q�x�(�`��;�V�����U�Z.����)�j)��\��I~����!������&Ub�r_+�Y����(�jÙ�9��9��h�`T�Q'ֳ��;��-�OGts����ޛ ݚ������t��!	�$l@.*�6(� �BDEL0�������[7Cݾ7�R�U^��X
j;&�hd0� *�DTEiA���3|�������o�o�=������~N���;�w�g=���4G���p���zsn8F�W��k��?�K(A��X�Y7t�L�=��O.������d�������Jg�@�T0�w�wO�Uy���������'��Ex�x0��d���K�����;��5��N�����e�s���>��W�bȓ����U��f��z����1��l

Q��I��@�Ș�$NA��~-�35�ǲ�����4�=X��]=#��X5'4��Ve�-��1WT�E�u�Y��H55�� (��/(�A��>P4V�Vf��#���ۻ�����\���F��3�)�ڎ)��Iyű�#_��fO^�A�7���V��؊��1l�]+|{���]5ƶ�b7�J����]߮&�����
�-E��*B�΢H;��f��#`r�z���������A�n��Ğ���G
l����,���:LT�Z�(�ۋ
���},�a��� '�,���9�sk��	 *��6M���gx	d?���}'Ha4�Co|��LD��r��,T�"� "�GU�fi[�E� f������e�Ls���-���w����.|��r,fgϻl��EH^\ೡ8�Af .+; ��gb�a�j��;M��	��K_�Ҳ8P������9���;4@�Ƚ ����<es�v-^z�$̆vk��\3������U�yl��O�y11�r���b��J�<�iO+*�z���7�,��t������j����z�"J�ű����ѽ�6�s,�@#[S{�^i:��À�.��%���/��0�j+2L���l���,lT;N�=��)@E�u��h�`L'�0��Ƈ�Fd���J�4�\L���	M��/���b�ӱ�=,��o�!� *���Y#�%5q%��Gi�RXr����q�(#ҙ����؏��t�2�r�P��"�ǋE�?�ma�f�/��S����l�rL�*�jM�j��J-s�$�4c�b���Y���ۄWV����䳞�����|�����:|�Cz@>,� A���Z�0P_�Aa"S�=+X�V
M�"��U*�c��(Tā��3)���p���8�m�'kH�����Z1�d��DӪt��չ`m��D�h�n#L���X�H��qW%�}����2OL�}���Mۅ�f|ޮ1n�c�b0�>_ބ BK��.+�ȍ?%~��$���c��Sё����4K�\�	�Z���s�8�M^�M��z1�o��V�	��	p�����s\{�E�
�D���at�&M}B���Q��R�L�{j.�A8͟���*��h�����q��Ak뭀�:?U�VWNs+jB�����<���p���8�`x7yP���v�+�+���EG�h�߻�S��.�t`���p�����k��%ӯ��������ӎ�;s�3�4md�����N ��ԩQ,zv�B4Mc���d�h��plB�9ǋ��mn���ow[��s\��"�[�h���X���7���T��N��b�SV�ct�)ɂ��ղ��(@�����\,f9���{k�P�z~֙�3tK\�g���6^�;}'�d�ۜA�~�`l����9��W���1��M{��z���]d��L2���� �)~�l�y�D;	���Eă�UV$�icU�h��u؉X�AԬv"?����HWAC�M������P��`�9��Ύ[*Mz�8��w�h6�S����6���ȏt��#���R�K�㱪��&B��$�c�H��`Z�k|��O?�я)����G�3���w��	�V���y�4���`�$�D_��ѧL
����3�!U\7.�f�H���q�F��lc"�4�-
�����n
8�4NI�.���~��F,��\�}&����U`:O���D:�;�09�w���Y<�ߐ+h�FY]��-����b�����ћ#�M����Fsթ�J�/�ˆ�A8�0d�Y�B�blN<��AxX&:Bt�Ȥ�qH�
����Y��o,�@��6�;��`:�cJa�6VQ��ɐ����n�v���X�j�B�	��� ��Ƞ�2ݽ��6�K^P�.�BȀ���n�i�;K��RMN�h��Z�g�i�7:22I�K��+_���=�cxG�Y_8��y��w�}�k���'�3�k!;@�P�\h>�}Ӂσ�%��q�]�V��'���:��3g�96���7G��PV����0l�P�����I�]疓8�aVI2X�ϱf:����0
B��;�u��7xn�3z\���H!4�j[e���.s��Y�=��7��Z}��L��|��2���e�l�{��a,�w�Z�?*���U�y-2��^���ٽ��,��DE���U���dY�}���s�}mҪ���~�g�h�|���F�#7�]6?�!@��_�C�r��aH��A �!�-��R�4|-ې�ؤ�L�0��(/�ى�2�'�^���5��/W#+si۲��0P������k�f�'I���Y:��/��0�����ogz�3����"���6�Ӆ	�&�&�D���03Q�N(��wm˽u>�6@������~� Nހ@�?�3?S�Ђ��L�:��� d@��K��<^I�\����F�K?DF������4e���]3ID��?����<��uו�c�E>`�@&������a��)� M���KS��nD���1��ʨ�9*�\Ͷ7�J�'�c*U ;6���������]>���-���(��,�j��ʢ#�Wņs�_���j$�E�μk؍�&�"X����*���1��ܓ�g˶�*}�_�2��q;w�t2�L7�dL��ݰ*�h[�\���X5��`a4"���P��K]LˮwP��E���F�(�(�^��-� ���_��.�i��o~sɠ���^f�M��Yo�vQ��v��?�M~��ʶQ�	�-�0�o��n���ډ�����X��)ҭ�R�@Ⱥ��!%; ��9�/� ����-E���5(;���=(�=���U�h��L0��Ô|�Ȕ夽h�_� ��hpb����#4��H��Ʋ�4Ҍ�=��@''<���U ��(���p=
azR�e�C��W���{��	c�	�z���9 ���E-�23
�N����N��R}+�Vy?*e���y,�	��[y�o4��&̱A<��
z�賙v~�'ծ���F{M�W.O{&�p����;G��_򒗔�#I���
��J�o4��{��.�S3��(�8N���R��a9��ن����k%�l<����`�C��횒2���?H�4�X-0���B�������B蘧V�� ��\�UuI8�įx�+J�Z��܃,6��sMl�fM��g�d��R�T���e��<�����i��-�뭴S��s��h0NW�;n�� .T_���<NQZ�M%�	������d����
c�;�!���U��&ev��?���k�gr�D<���7���\���f����na�<�ϻ�գ�������6����A<&� �Ǥ�Y�E�E6�Y8�M�����"G5fA���Y&�M�RF�)�c��(:�ع��}�|o�">�o� ������S�f�c�MԨ�>��h��r��-S0�{���)LxV�k����*�u�ݍ�zt �T��P�l�"4B�����<k��,B8kxʼzD�CN�ݝ׻ݽL�2���T���.�%]qFB�餃���R�jgdڻ�}����{������S%�����{
�#�����׷��嶟7'����v���+��~�n���"�����#$U�4���Ѱ���D���0���|�)�L�wz�H��KAݠ �j��5@q��F3�<�U��V������=�3�B��I&�B4lL���BK��6i �}S��i�0s�e>����~�b�G�^Ď�G,�� 1�Fަ��o�����^]�e��n��]�J�C�)@e����O��v�Q��ʫGgPro+�$�ێ��(�S�;.��i��e-{��8�����O�Y��/�՞k��2�D3��&v����,��A���pVPf�}��ש�h��qg��eV�jw�I!��f�x�W:��\h��wF,��E�y�����6��5�<��ܡ���%h�nLR��c�U#\���>��	��w�q�c�&�c*g��>Xm����J�i�I;��"4���ͫKt�g>�?�9�
ܜ��e`�D0�v>����ʕ��_��W��=n��꫋�x\Rs�tG�F��%]W�㤌M���z@��5�J�c�C�6��s�E�{Ht��̅ӱ��@�z�T��m�ud��, q^���] 8�{��ģ�a������ݑ]8D��v��6-+#ۅ����e/+�e����E%���!J���[M���S��a�G�Z���1�����\��SI�Y��-����	S�b�5��}a�6Cm�G=��%n���G�:�!�>(�/B�L94ˊ�	"���H���/.i�=&>uEA�T�'F�X�D����b��B���b��R���ksE�zҧ��ʦ��k�v^�7mf��QL��;�%师L�]O&�1� [�Y���A|�pD�����^�c�
�y�!� ��Q(���zU�D�Tl$s��0)�.L��Fq��F1�,N$?�W���V�>چ�=���1�R$��}��G�?�%������kvw� te�\�3Ep"����q�dh��"�R�[��L
%�9�)��r�������X�7��=>򑏔�,jU���U�z���/�ʖH�Kq���:k.B�ƐH �U��y��[� ��S�{��Jb-�=f��� $*��|Ϝ�t���"!� cY+�ۨ@��A|F���r<s�v�2]��y�5��(ؤ����,��M�Bc��_����D*f�c���e)Y�� %� SBa�[@����枤]�<�?�pݤc��6Gee�N��-%yb�D��続�?���.� 0B�,��at����A ����P'&�c�Q\����F3MWۙ�<M![hCU]�]�N�z��C0k�f5�bW���/m}�������B)l�SC����S�0�R�[)��ַ���[��"8���7�s$Z���b^q-�^��W4��?���LJ-�Ë\��o�!��;���M<>�������Y�/��/ԙ6�����ۿ�|�h �gĉfv-u"xVk##{�~]�X����h���g���ݐNw�D�`�@�q|ڝ��I+���Bx@�Q���&�s�O�6��qkY]>��/��-x8:,��
F��3�nR�v�D��M���6��Yp�O�QR�J�!C_L�>���ժ��n.�.�D����t%W}��R�Hdz�k��R�?�)�cjB9���5���(��Nt��f�|��8�����qJY��y��h�F"���\�hv@����|���)�!�)"Rw�ܛ>@���2������E�z�օ����	��Dv�!�耢s#T�5`���?C�l�Q��R	E�ⲫRЮ(%�u��Xcu����&HT%��4�cݞ����!H�ņ�I��G��o��b��ZT]���<P�5�3U9=��t|����"��v^��MӁ�c��^���)8�n��v>� S-t�o���`3��cR�}
��Qȝ!8�H�x�32�4��_CHQ�-t�-���)�W�)�ۍJ��`����h�����o�뻾��0i�*h8ܨ��%s��ұ�9}�s#G �`)���	�J<2�_���Q.����uD.��)��;�wW��JO�����>����ǉ��|i0O�J���5�#��]��0��~闦�`Z0^���A]�� ~ғ�����e�����#�fy�Y�e����<���y�9�	y�Ь~��T��\����'��K�~J6��o,��Ŝ�0��O����
#��bYF�ٽ�mo+�F��s 4�!,�� &:	r;M�鼭�$�W����q�")ʠt"" _f�������E����W�(R(sM^,PԞ�gʫ4:N.��$q�M�m;�:4LIU��ϕ���;褁�(��Ƴ	��0M���5�3�-��=�N�qڮ.��㦋�?���q��(h��;�EW"*�~���A�|��v;,�55ZH�� "~V�[{49��
A�����s�"D�%�a�-��=�g��X� j�̡4�%R�G
մ'_u1��1���_�j�T?P�	j�g�.���!Wڬ��a���bǪf�}t_�e������A����Ԁ&6e&�d���:�B4�ݗ��<Um���&�r5)�Paw��8�.K�b�l%�ˍ&2�Ӆ#�\��ϟ}��jW�h\J�w�!j[$ktk����O��X�+�fP��v��-��l��KA C��^��-37,b�KI_L��]�W��2�%��Ō�v�d�vv��������B=A���v�"h� �xf[iFМ��]��,@�%§>gdM�}ҡ��X�tGw�#g��hj0�]5��l��kj�I�Ţ�1��y�����h�B�`8�ť,����K���N쬧��s"c`u��(��03���:�����/�1<NT�����~�4�t5W%�ۧ�}�E�9zs���7��|)�0i����Jngb�_���6���Rt�]�4ϔ��|'�~���(��b/���rG���6�4a�Ӟ�'�iF�(�t �����^�"��xv���6k�'�%Q���ފ��޽9��"�Xf)�NR��;�	���g�-�� ]�,5̀�&��6;S�+�)�y�ܺ��i���,9�ߏ�v���*�j&�E[�_��[�id�k
_��)��T�S0�7?�"\�s4�n����s��m�o�t%"�p"Z�1�t%��e�>Ʌ� ��h�Vi�Җ���b�j�U#�e���J���,�(9���P�}��"T���lQ�z��E��������4�=}�������v�&2�kߏ)[��L6��!��<��|�WVS�f�-Qs��t�mH�q�/�ڶ3^W3�Ϻh�̣4�@�5_��OZ,�WT)n��q�6�>&�?*�i< �_j�[���ߙ5��VЋ��൬qꠤ�@�D4mx/�;Zd��g��8��g��Y���^S�Y?�(��e�Mڹ4٤-�g�g��يI�?���z��皕U���lm����W����LP�p,�{�>����e։��&e[D0�(������E��ϑ߉^�l��\�����Tצ��Od%�QH;o�
��i�NԘť<5/�R0j�����z{�4Zx=3�fQ �u|'�)��I>���=����{Q~���_.^8#{T���vA�H�[��Wzڋ�9e��B�n�p��z�R
�X(���T-j�!c�ex�� ��n�ݐ�\]�1�M2�� ��|�'���>��ƿm�!��iCS�7�s��u?���S8���A�/��E�6u2ʇ�s�ZX���m�hš���W�Q�G5n���J��r��v{啋���>S�]���9n�	B���N2R��%:�{��˩ۚ�L�C�Q^�k������	`��5���;���9g�f���U)s��Hj��>9��h08}�Hx8,����7L����[ؘ�v�^Yo��<;����J�ꖅ�U?\��xu:"�.Ls�/��m��-J�W`��9	jЫ<��|�(�A��\��������&k�f��j��j�,sRM�A��XMl+��^iphǃ�����N����ś����]^@�����~l,P��]�{������X�
9�,�(���@�xU���Җ��+?�b��Zjx)�Ҷ�ɝB@��e&��Ț���r#%��!�Ŧ(�y��ㇿ/���K�M��a)ۂ�^q�Q�#VVze��7��;U���W}�_o�k;��&ج�.i���$ۇL��C.0,F��6��w�@�E��*`S��d*�tl'����v�ʩ��DE
�p�B@�L�oE6�(�>�������!(0 �ͧ��\�Y⹇��t۰�V~����?�R�����0��֊ݝ�V����F�=��U� �[�M�sͥL���!��妗YQ�1��4�ɳ�δv�e�	XD5*�-j�^���IJ��m�Z�M>��q0o���0m�|��q�k�igتQ�>���"?i����]r	\S�%t����n��6���\!|������ŧ�����`�ln��'ڎm;���}�U͉S��yV��<�9�f�<t.e�O�5m�LΧCefW>�w����&�H�"�v���
X3�,b�03���J�n�"�SX/r�uۇ��b���R�+>��`d�Y2Q����.D�`/��������+��x��;K��,��u��w��޻]�A���ܫ���-2�a�p��=�����j+�vn�N4���#�B�����Љ>3�_��9���=c��
�=��%: �(�+�T@��m���C~OM��E�lw�-��kB���q�N�癙�TP�w�#Jfo��������������<��>�*(mY�X0�w��m�7ƍl��6�Q�_��<�1k�[t<<� _8Q�	a����.#(`�,jz�K�j߻�xgb�U��	��YE�Gu&��QϘB*2}
&'N2,��
��#���
T�B�.
]�*��Q��1��S��~�{��ez��B.l/%R�kʊ�ET���b۝h1�Z}p~��Э�쵼�}��f�s�����M�$x~����Ѣ�m&H�]p7N5�'O7ۣ����[��k>��ϵ���| \��=6��x��V���Xi�<��$66P�q�P"N����3�{�
�ź��l��`'�� IW�RX�9���k��e��A�Tf��o���ϥ�'���Ԗ��0s��6��ŏc�1���񿌜?��~��T�a�i�>��n��{p�w~k\�z��fY�9|�ӓݖ�'.�6P��qX���2��}m)pMiL�����z���m�D�aJ��d*���믟�.�`��&U�e�d:J���aS4��ך�]a;&&��|��3,C�&�'��?���/E�a������l�����Ye>� �F�w�£��o�Fi�y�9gx��XG��h�;c4ǳ=�Y�5�}̣���<Ӝ���f������|��vY�G���k����<�-��ۅ���͕ts~�b���{��8�΢a�x��#�wߗ��Z��@�0ο����h��O�Q����UĘ����}�X5����$+d���2������ȗ*f�����t�97�'�!��[��N�;0��^(��s�1��1�L~��~m��5�����/x��_��_�.|o��Tx��	��w(�A.���XC���:����$�7 �Iz�t�R�m���fj��n��mM����*���vyQ���(�/�R��~��`wh�ߩJa:����#�!9��� 08���9�( �+Ì8a�hv೓���A@�L��炥���h#��>����	R�fҊ��x�ϳe�	߻ןU��M��`� Y_�Ew�B�h�h�qeԎI�]�Ϸm�Ex�9��;����~�X�&�/-/��yT�4W�n5""�'�����>����~\�ܱ}�U�K�PD?#���'~�B9�w���uP��)���.�C�]6~jc���F�}���@Q�����f��1i�E�r'�e��|�3�Yd�;����ۿ���w�/�����R_�
6�Q��� y�<�AQ�S��]�R�����q-�sG�]I��+��3�	l������U$��oM
2��ЎRhhc���F�S:�� ��R�w����=�!�(�e�e��e�P�Iv%��%�禭++Q�7���P6h�E��̕i�Y�U��Z��2��6hW��z�3�'×�3ĉ��]sU���'�5�|Xkm[��^iE�U����볛줟v������jy�-kZ����Ҿ�a1b<W[�^8-�w`E�h��t>��4U�4�i6s.��N��hU��ڝN;�N!�b������W'sn�OĶ��&�;��ֺ���3"@���}��1���d$��Hǝ���h~q~z_��fJ�6#Tv��H�3��#O[n[�>̰���ꇚ��E��Uk̼�J� )&2���k�����!|Q�0=`�0�	"�2���_�I��P�.yL�<2�q�m��O鑌b�8�hXz�N����.���ҟ8i'כ>߰��J�ƈ05�o���$��L�a	^[��V���7�9�(o��֬�֊ѡ]^�Ai'�N�R�BL���s����"�ü�ͻw��-z�}7���X?�A��&�Ź�%��g47�tS�� &���1̽Պ]8�؇i��|�L��ҾX����eqWO6����9���
��z�)�^�$�r���s��PG� _lS\��VɬF%Cw1�/��y�<k����x�.�K{�I��Ьg�eJ�O
�����c43�tǉ�@Л��p,C�G�yI�W���N�a˞8��Rk�j��o����kMo@��N9��|�R
�Y<Q/�)h��Z�5�ݳ�"_��˜�ۜ'���e���_��c��� bh��ԴhLp�y�F���%K�*�5A�#�Y=��w@���	�ֶi騿���J8��r����)��N�C�U���i��A�a�����a�bl�f�m������l���`L�搮����Yh �LM�PD����:��eֽ�����i���f֯{df9h��[e��qZ��>�Zi�ޤ��j:����M����iX5ū5u�y쬿��,�t��� ��E/zQ�z	���# eK���ۈ�S����V�7��SKT �N��W����	���m��6ڝ�{mD�x�4U/8�g���C��ԙ75z� ^�4�{U�/�t�0�N�����jd�Up�Z�}���,4=��௙d����H��5tI�x��X}�.ҽ&�����V�)O�����D�p��¼ԗh�3�r~����y��^�ۼEt���K�*H�-5�8�)�&M	_�5_Ӽ��/-�  b^D��	�_����#������n��פ?'�(iZ��Fo�=�Ӗ{��c����	��1.�	Qgޘ.;�Q����ˈ�!�9Z����f����P�e4O��b�Y���N�E(��e�E��^`�۾���wfo�%�gԢ��T�����7,/2��ʫ!ss�����lM�d�]d��Z4��T�zQ��w�~�Z�C�JS�֏��-�B����w��(ur��~���9S��h�ܹP�����g��&�ű<L�+�}���s7����(-3�߆�X�^��f���?�8�D�؀�|��ߘ#>��UE�'g�X������y��"J�j}�A�<�;o�^��R#�"�g&�C��{�S�ؤ05[n����1KfX�p�����^��V����������fH�ۨ���K�,1�O�� ϲ)׿մ/Mf����z�����"��:l�K�/1�8�	�\��FL�<�D��g����6�/J�Ub��Od�>ZieоW��!j[#�sDz�w� �{P���}u���N�'RP�@)<�	OxBY�f�5�H�
Z,Ę��؂Q-�jA�`�+���v�SK����M��,;aݧyݬv������f\%m�B[��vnvz�6��IXk��m��ˠ�v|G؁����Aqᵂ�x��乊�btI��y�z�f�f�2�s�WW�ټs�^��j��"g�aH�W�V�ٝ�цMK�j��Y�7?ב^�-A_��P;X_/��hF��[��k�hgP�K]����n��������N�ґ����<xE?�яN�T���h��l v�uQY�}��t�����p��k���.2o� �>�'>��0YM���MR=i�Y��@0"ǳ �����$b��}�q��CaWs��ZG۹^��ELX&NТ崇�w���������4=ܭ3������I2�,�h֦��JU��n=��K������,B����nF�ԞX/μ��|s)Q-h�����^�ѵ�^;�D˰Ay��C�E����HL�ٝ!�y�i�R ��[��LQ�ݐ�=$V�v��;"H�'Z(�Ȑ��t�{lF8��7��M���}�ו�A��[��ɟ��TF�j�L�x5S�
]�ߝ�Y���`YQmy5ҬA��"��m_���<ٮ<��q��k�d3ȇ�F�j���|utD��f�H��2��!� S:�2�54�/"S�3�;�b�
�4�X��A�ٸ�����r-�d�Qf%���j2EڊP�Ǆ�/h/��xle,Rz�y7>۾6������2,}ɤ�=��Q]����λJ�Й��������R:mP��JɐM"ن�D1F�8���x` o�dʵ-/�E>W�n?���<ِ�����U^Ÿ�Y���"���k����M�y�{
����y��)r2[sY�h�\��0��3��̴�+�%1�+��υެIgh����xf��E�u�����2��H) $m�ޟ��N]ն_HЗ�X����3( �e�����j�S@%��]]�(+�)���+2��+M>H2]�\|�������䋿��(G�xP(�Zv���(p���I]�9 ��5r G+�Y�r7[&�s����X��s]�|��y�4���l{d�=���n}�G��eә�w˜.E��Z�{w��8q� tn�m��z���N��7�����Qn�4��(�jd�����V��O�������wi��t�V�V�B���|+�g55���u(HL1���� \��1V�Ԅh�*yV��!�3Y["͌������z�)/إb	��h��}�@�� ���y�\uQ}�D��!�.�q�K�Ej3i2��)��W�H�5���T@)� �m�D�(�G[M����N��_��_++*�"H� k�9�yN�Mj���R͟g���Y����Ⓕ�tY�&pPUwl{�^�k��.��R�rR��<�h��dz�5�p���_�+�n=�]���¤��2<�2�^,'Ka����8�����]dW6�;eLh\Vxe|͉íe�r�������M�Hr�X�9��7x������-:͚�FiG�R4�9e��B�ڿ��碑%S}>�Mm�9#R��ѥ�ڛ���"�5�P��ڃ %�־2?WP.H�P�P�Unh�Ȩ�Lh�����G���##��X��j�LS�A�DW�0�Z��&U�\� V>�T���&��*`�O��OM;S��E g�@D���m��Y��L&�h�{�*��".�q�r��$�x�h)LHg��c�J�QSH:I�N.�9�]h{��Y��[��!@���9�i���}�k]�jd|pE��q���cĿ3�)��z�_x�QmW;�+�Π�#��X�{���1�P�k֡�"��p�:s̶["��t5{h*��꼁rA�9D�]���	��^����������� P[��L���vhb��n��g�1���[�ȹ�};�~�GG,�'�������1v���f��Pm�H�,�a�h��a����ud�h��1g�2I��b���� ��i���\]s���Y�G���+�ղ�}:gr��{:F]XH(H�
�<�����a_om�0���ń��.D�����N�s4A�͸�Ψ��Y)���NwS.qÍN`�ž��#�7�C$/U��1�Ij�R�Q�m*D)e��X���s�\�e���^���ҧ /��9�����b߅�g�,�Bʸr�����e1b�	J��T#��o�ʚ	�j9������ZDN�;�>M��Gp��ϊs枳�����!'u2\��$(䤭O(��iO{ZA��z���+��+eP�v�����"��,]�=;�P��D�P)�Dz����<GT�0�ڳ��(;M	N��;�6gU,��ue�e��_
���{��p~���Z|�GeM�h�����[�IGc�:�.�}څ}�Ef��˽
���/e�ܔ��r�M;����B�6��p�N�.�s-CN�Ye{�.��{��N�E�<��gKg|���[%��p��/������r�Y���H$#"DЖ��<��!yuTJ��4�j���R�M�x�����4L롧�*Q�<���D߭˩
��4C;\]DPt\����o
9��5�)�'���Q,ЬP��j��^D�z��hK�p4�v-��
�I�v��L�k���Q;B��H���P��
�,l�ئF�t�jt�n�����-���&��m���λ2�<2�t��h��>z&5��?�-�A���d�	�V�����p�Slė2�����^�M>5N�hj��0�\�S8v	QH�r>A�O��(��U(�춋߻ڂ%����8��TL�:|F;��>�k��v>EE�ڴ���9� ��s��B�y��_�d����V%Ul/͸�֢sk��O5�U<U�o{�ۊ�Fx;6=�ڗ��t��b��	�����g���:���~I���T��ez�#QWmk��� �h�n�����=�jh��`l<�d�L�kT�.x�q�[���k������@a-�^�p8�y��F��C�u,뱆R t
�м�R�L�ؕ�=�G�]>��8�H�D��x�͋_���)OyJq�s?�I�"��L:�dSon���<LԿ������s�S[8u@�fd����P"Vn�=�F����Fꕖ�~��)�)[���
_h?��yt���4N�m���w&;p7:�,ҥ,όZ����[�����y Ӽ���E�%�XcзU��ַ�=X���B@S_BP!�U�.k�祶�5 ��4y֣������R�ⶻok>��6w������Ul>�'٬�Ϫ�:�h�����I5�T�ۢ�v9��J��$����E�y�7)��w���σ}�t5J�t�u����O� �2���1�"{��V�yx�m�]4��}i��j�Ӷ�誨IS'*�*1�S(���^�2J�b~.��Y��B\M��y�Zi��4£�e��Y����2�Nc��[�~6��vK�ܼ�&�M��_p�K�q9�aA�<��z]A�~�|
[Mځ1I�����S����e�i�ά`���#��hsí�R�l�����D8����T���p�ݦ�Xt��6v�N �ź���ric,���܅�b�OA�^�+��f�ʌ���[o4�s�pυ�.�t,�5^|-q�r��dw�@�Z���!�4h##������y������<� ϸ���7*��iW��v��}���-��<��YIw��������OpW�e�?,]�4)�>�É����5��񽴷�����l�w����d��y�(��D���0��Q[v���0��cȘk��m���a��/'�?Zj�Xf�Q���X?Lx0KlV��A���Mx4)��Oa8�3�F��E,8�i�o���qͯ��U�ƌU��+
�Ġ�@9bA۠��ݬ���e�_:�2���zj�I��7��w���dS�f����]F��r�ڬ�+�n�E+Ee�V]Z�;�����-ȳ��kHa�M9ߧ��Aa|�tX��7��㘳��ڂ35�cY��ΰ>� �L��GQ�0��u�	K�LQ�暃N��)�ks��ze:m쾬��ԟ\�ܹ#�,cc?!��(6b=ތ	������'��~�p����3��#��a�'�2S���2� ʪ���'�����[D�c�"[^#�-b5��a͸�	#�<��7M8˦��	SE�Wb�.�8 ����/~�#�����N�$�R�	 �;�9䠂q�����A:
JA��m��2�明<K�@"E�נ�eg�Y�59�FK�#.'��z��)#Q"�6�E��2�3ge���A��I�>�@��d�Q��F³4;�`���s�w\����1��e:�h� �}�0�=Z
s�tJ֛H�|�s҃t_P��*!@��=�n�iɐZ��Y��g8��i�.{!��D�ڈ�,6ߥԤY8�����R����Z$�����dĒ����^��xt�s�q9�"a8�zT�.C�VĂ��fM��`�ti�|�++�e�4=d�nskqw��A��Lz����.{$�l�3��(���YK�e�N]�X�=��=H� ��-k��)3T�4�oC�F mpt��� �G���W����]֮XF2��8m�҃t�R]WSD�,�G��eM�4A̪i�`��^��0dQlw� �(�y�Ö���j5~�#�K��N�3�򸖉%x��u7ǝw
O�@O��-�Q1�1�n��*b�Z�Z,��?큦�&:�Tt%vͦ&+�s���O�B�X���7E��	kvXa�ο�[.����g=�\볟�ly���}��ԧ�xn§���չ��Zͼ~��G���_��e�6�~��X�Q'+�j}A����ig��ǔ�F�pj���Ju2�	[1�0�e]����u���S@]A�߅��~���wwW�L�L��N��v��`K��
���3
����������˱0E���暹����~��C�^L�����^َ�Ҝ#c~��/��	QGR�H���]OO'�&]����~i/�X��)�ԏ|�#�lN8ⴟ���6Ox���}�c�w~s�F������2&��{�W���r_V6d�~�~�,z*�]�X�RO��E���GuD@�-vM4�Lهf�AY;���4#~��`,��a����yO���l/�.6|����y�K_zA�^H��w��쀮V�M��Me�,��q�-6�u�u��L1���C<:�I��")�f 	1��l�����&�Գ�W�Y<\�Gx���!L�!��gU~h�������w�5KU��qYr�@(���-8��)w�6�ߝ�3��c���*Z���,��g��1���?��JSR]�oY�.�ܭ7�??/"3��_7��><�a�5��nj����<7�����٘<�n-��b��\lsOC��eȚg���u��a�������i�^���ovmI�0*C��=���뻦��D�	  ��8��H$��=*r?����]�2!�dr��
=�e��d`�8N
�Da�f���@��x+jy}���+�Nn��/����_�����Yί$c�	'��.�ۏ��$"�V0��\Y�hrh�ews�r�pr��Yu�_}��g?{�N���N�c*J�T����+['���~�Y�A`$�U[��� wa�w�Ff�~��8��b�
(�͢e��V��q8�D��s?�Ð��>5:$N����~N��W�m�|ge=?���^J����C�9����sKV���r3�.�F"}�e�p����	z���wP�{�s]l�hkɷ���P�U�Ml���]��1���D�����`��,b���P�P��-����?��He����-������� ew
8(��JN�܄�3��}��Y^�.H���18�D��#%���z��D�j	)DT�sgm�:n�Fѹ�0��6z>�0�dͣY}4K��f�Ft	�d|<^j�ٮ�C~ss^(5�	G����l����D���D�:��oc��un^+�v��[d�耓���2�L�JS���c-]{g��9T�at��ǧ�`2!�q�bR}��xGE6��N[0�0�Cާ����� Ƴ�Șŏ������|���k�A�v�5�R��9�g�g�3������|ڥc��>�f���O���J��K� �3�Ф �G<��g����~y������s�|����s Pu��ϴ�g���s_Y�v�絉ľR�+�E��F�h�j�-��OԶ�h3��^��q|VD�����s��ۜ�v����{,�Q�1���p����&,RϫW\d΅�E^�d���;��LD*L}򓟜��yԤ�K`1�;����z�.!Z��mևN{���	C "PR��!Pm_��W�sElLZ"@wD8�������"-=����W
�T�^� �DB�ig�G��ɾ�Mܗ��?��?�jg�+�Ȫd�k�����;���R�3�#�+���s�M<�O��2%�c��3f�A�"���[�G�Q���f~�nL�ᗾ���f�����h�pck4?ad⛕f�4���V��±ߞ3��KkG�o��x߰��h&;4􇹡�{뎏N�=�sVBp�"Wk�뮛2h���e3�*C��V����t�pkC21�a��z]�r�Z������Y�&K:��	�E�$t�-�w��%��g�4!dZ���6B�2?��?X���C�6M�lV�cr���?��?l���7��G����YD�=�=9��p�'=�I�����s�."Q���o>m��2�|��6R�xj��4��~��ӟ���ܐX53B4q�9:�k^�{���d����VB��dK������*��3�)Z�&�vv�K�0G.t�~^u�aj�ӄݖmͧ;"��+�&4
�f�����q��^�"������+8e�D�V����Hr?<&2��C�MU��J��Q_;횵�Lov���I�9G�� v�/b|��V��ޞ��t��6����
=�^���1��z�0��8`���3M��D"8�ːp�gد�_;�Db����өC�E�w����ɟ,h�6s���H�tJf	J�r�]�j���U;K�gJ>�\�w�jG���(�:�Mb)Fnm3i\iZ�MEq+x�F�oƂ����u��|��R��C����=�Π�*���_U�z���j!�9�"a�y��;0�,A9w��x]�Ʋ{�Tx�|f�i�4�B��n���&��ϴ��c�� �ڎS����и��+
ә7c7�CS-���&���h$�h�UՇ�8���Y6��]��[��NmNgf�ʛ��ߜW��g	��P�	߳�9:�ϋ�!�	�~�}�N��p�}�!P��ឳ�!d��9�<���u2���
M�sʕhmV�LI�W�0��=o� �����<T� h@���f���:B2p��`QbrY�6�Q�i�L�,�I_�r{�e�i)HLڊ53d���g�`���r���§�6y�g�������l�;�<��7������ʃ5�p�#�򾦨�M�}.�5_�}s���t($� �Q��v��W�:���2Hw8����>lrw�r���� �������nj��,A��9�\���Q��ʛ%���.�!�������jXm���ѿ�g��o����x9l��`9���:�>�Ut��G�gݍ��{N��B�{�Y���i.��I;n�B�Tq_]��}�B�b��3u�^�1�Ye�� �\S;�o��1�����Jm�>��}p�f���N`ϟB.c����p�ĩ��#8���ۮX�G��_��E�m��0���Ɵ'N���:El�z��C�[�Wځ���������O�o6��@H�
(��#���^��gQ
�d�4C̚��T#s���F3��,L��U֪?����xS0�M�߬�����57�!f<�QR��]���&���|� �@�X0��(���-.�i�2t�"K���Zf�5������E?��,�̉y�y��xl�.:(�Nw���vk��lU�MlX��c���5�=(��{?�o�3�><�.`��x`,�/���åJW�g0�H�K�Q`��[����x�rY%+�O�i��N�ɬ����s-��~��2J4m4��`GmT@&�M�B�&�	�̊�j�p1�q��fۛ��\��!�+�k��7��}Ώ��E��������?��D�T�Jy���W6����y �v�)�3��1�:��@�_5�4�0�,X����J�����(�r9
�Y�9☣#���(Q��nc����u�f���$���Ex�&��oW-|j�ϴUVz�?��&4�I57S}s�s��~��e"�ݿ�w2�5g{2 >C�2LG�Fĵ��ZLG�舮j�D��h~�F������ʢ`C ���O�8y.���^N4eg��Z�ǋv��s�S�h?�<J�-��<��գ���?���������FG(|�9���Q���-K)�چY��5A�)B��gj��>Ke2�Dg ���K^��/3�Ĩi�)myQ'"lGC�	�"���U����F�������Yk%iq���-�poT�-�r���������=G�f|h���8�d�X`l^��;�SJ��=7=���f��ZAo�ۋ�&��	��-T�^�{Eo����/=�
*l�L�.{�#p� ߯��B2<�'|*�ʈ�&�Z������o.P��Ԝ�����e�b0N�������O���t�!h�P�i���<�'ٿ��d�x�[���t�ME b>��k�����k^���6�Z�֋�NJy�y@FZ�}����T�1��L�X(k�A�_�ѧ�7���T����˄�t@�2�|�䳎tqBԦBvT�cy���٪� �^�R0#����� �ڼ�v`OA1��>���
C:og06?�W�5~�}�v��?���bC����N�-�$�����P:�r¨T�m�p��۾��u�ٜ�F��o,�h�(�XC��y2����V$l�En�äE��2�H��C�d5�ְ*kB���>�<J3�Q�}`yO�^�	���-��@�@���f����@\s� �T匚�|4�v.�y�.�4M[9����7�&��O��V۝ʱ���s�����#�A �!ad�=Z-6�V5;�z�[� ��I������pТޖ����j����V���V�A�c#p�fפq]�`bׅ��i�Ө�=+M
�����h��*��I��@��G�o��h&���� kRNM@������M�]ǂ�W�����i��N2�j�Ь�DTƣZx��07�
c���|hz���}��i���f����]��a�ɲ8g�	G���?��X^�A���w|�\B�R�m�s��yF��3���:W������3�Z���w  ���,��u�ˌIx����#�mv�X���j��;=�\r�
���b�f�����l�����6����VVWoﭮ���6ۡ���������p������m��j��+��S뽕��5���i�;;��#�7 `�A2��	�l2���5&�G�T_p���*�I
��x�_}\�cQQ��X�t�+���ɿsҙ��9 :P��j�E�u�tMYD����O|b�7�aϹN^�Wۍk[�~��㢌 A00��ء�i|;�n���	������_�*~��#�_d��\� 7�P����r�"�f�X��v1R�b6�Y[3W����Dۘ��&5P�
f}]�އ�%��9��bѝ�H�`^�"��k�g��m�k'��ub����S:<q��m��S_X;ٿc��~��Be{pb�3ē����G�Νy����Sw67?�<zg�������U�Q���';E��q`Pj;Q�l)���t]A1KT����S���*t��,�嗿��͓����0|�[�ZTP.�T�W��_J��I&���,2�yf�!ϯ���'��֎Ό�p1L4g�jީ�6ե��%��Ї�Ї
o��u�+� t��c������O�g�9E�:K�G{Ws�}���'���?}"��'��yâN^��m���  G�\��d�A�ӋBY��P�m=6�����@x�I�Y���w������^�������m���W=䃽S��sW��~����}��Woͺ��7�w��ӟ�X���U���Ǐ���g�~v�̝�\��~�a�!�ع��g�_��Q�dK��yلt�#DE�:�p�Y4H{h�MoFmReco.���;<ݿ�˿\�b��>�,�js����p��F�^R��tX^"�e����?۔��*o�ڋ�~�2��~����0}I\�/��/�=E��vJ��K4~�߂��|�0��
Jx7��E�6��p�s���31Ͼ�[��h� b��)��
��=�s'�o��oO�AF�dx�qҡf1afTI�o��!����k[�'O~~p�C>�y�U�>����g7��I7��|F�י����������?_������o�>�՝�����>��1��Xg�G]�&�A�ƫ��1�9�����_}��W��`l����jm.�����8���>�,�(��o3Ѳ�/�2����p���z�긓>���x�R���ߘ�@r� �qcƯ��l���4f��� �g]5�״�BڬYl�M!���E�"�se֣ a����0��PW�Im��� ��"��	��`Yσ8�<Nx�<�茘Ҟ���<-C�O4�VV7�n���֕y��UyO�a���O���es@������z�?񾇝�����'���yp��ן}�7��5ɬ+�dҍ+�MPڴ�İ��F+Ӻ0�[Y��U���:����Jʤ�;���
�Y�9�<8XP�x�ɬ�ʻ�L8�u/�^���$����\}C��&�B���{�)��Vp���l�"{�bV`)���ؤ&/���3��50�]_d�K��e�R�y�o�PTô��8����!g�S�z�э�ŝPCR�+�^XD��1�e����>���2��S�G�	���˦�&G�.K��y���P[��h�����8��s��݃��������}��s����?�����So��/6���hV������+7��*4h���v5�W���_�����f=,��$ʢ�g�����ZA��ŋ1�:��Q��D�:��^&m$��«�C���6���Ѱ[!L�v�N��2R𤗹F���Y!j�'_���8��Ƣk{l�7Qp-��]��y����1HMH�X��6�d��BH�b%������)�B��O��O�1�
J'S�^)�f����q|�jkj3�A��f�5zh?!`�ۍ �������<K�]����C�e6`nQ ��^.�z�<c��9�6:"i4���������t�ݜ�m�������_y���C?��׿��8�������/~�CkW>���F�ίYkzW�{L�Qz;�����~��8Iz��W�cw���ʇ4ḁ��l'[����؛`2P,�N�y�BF#��UY'�s��ܢz"��&�\��
�+��d.��ȝlf��f	���RsrմL��2��3/{>��
%��k�~��R�ÏV���L����/�2 �dLX�+^���~�Ǧ��2痾���ق�O_�QD�=��y�5Ρ��,��c΢��B�9��w�wO��C.�5�����/�����i�maԻ��	���l������s-�:u⏆W�~���'��/nx���1�-?��}�i�����`�����\��5�vm�[/��j�;�bP�K,�����|Q�e�7n1L�BH�Gm�fM��h�+91����w�|�+���+���#g��.θ��L�]"��Х.d�Ѭ����P-������\HDU�%�	K�"��^\􋠂� 8ٺԾP�����7�\�ז�(��HQkk�ׄ�y���β��"a�-����x�k^S�jS�AHsJ�f@栵34��X���Q��Gl.���j�_Yk�������[}�G�u������1�����������7���w�����7�|F�>ͥCc9ܯ&�pƼZm;��xFab:�TH�1kJ��^W	[�{v6ÄX�l�|�:"s� ʁ	ͱ�`�~��KFcEO[�ahV�X~���c���}�s*���lbR�Ǽkxy��	� ��Ř�)a&~�@��)'��3Q">����j��BV�<@˃�A�%��>�N�����%�A�_���xz5D��i7f2i������훠�᱙#�Q��0Zoz�'ϵ�����?������>��+��k����:�I+۫덆'��z�qt�Q�+��F�J֞� �|�b	�1Y��v�%]�|9k������N�L`������L{��f��]:K4��%P갠K�RŮ�(tXD��<s-�<A���sSP��=Hm��P/Y����wY�s��� m2>�!�KPt�9�O�������p���f��F�)Q�O��@^KM�P66���_���1�>�~�0�ߏ��Go-�-�ڇ��F<�/����=�~ss��7���'����GW��9�[��~�~e�k�hX�hkL� յpxY=M䒔�c t�������EH'w�5��
��|
g�.*�Ӗ�m���1�����.aH�h��P����&lȖ5��:�vQ�)L��&<���}Qɩ����6�%@�
�.��������9>��@����m�s�B����z"�Ed��@ �`$�>,�98��>ۇ��h%�$�����տ�Վ��3X?�?6O�x�'������>��kk�>}�7�����`篍��2
+X�{��E{J��1q6YMlĮ=o+�&ֶ�M���%9X
\���SebtCdtr-�I2�L]�EyH��ѱ�%��`wCxX0x.P�QT����R���j�zm�?�Y%���+�.�c�V,ͺ�ـ���O�I�L� R����wO�]��귄���h��)�G�`d��،E�HF�:7Zլ���|��˽<f�7,2����}��U4e����Y�F�n����룍Sw�_����ɵ?k�c���_���'�|���A���͠z�'���kE��}�c�⢎i }� ����sY��\�A�;�
VO��vf�>�/�o�����ȝ!pȩ*v���\��Q�}XA</�������2+�������&������"�1%���a��ʐ.$D�5Gl�'�$�߬{��?&�5�a�8�ۺ
A`E3�&!��I�hl��qaX��25�,�!�b�@x��n;�����`XP01^�G��&t�q�c���� ������\u��'�z�؂��7���a}�����m��k�VUMV��N769�C$���K���-T���:Hǂ81�����b���$�)�c�Q�Ҹ��yWgse�a�ߨ�˖1u��lzk���IO�hٰ�>�$Fp{\?�2�5�@�'Nxۤ����!?NJ�������ctpZ�ŅqY���^��F0�k8�ue�H�X��E��'�s1,cK袻m��rA�]D����������_�k��5�3]Y7��a�f��7h@�]�ɺ�j���?������X�MVȲx"��{��8������Bxp�Lo��.�������k����$e��++��N�E��~oog��a�h0��������V ����1eƆ�X�(D�M[��ݔS-�z7[B�s3�;2�B��Y���jS���߳��]��\ՙ��q h�:�U;v5Na�=�+�<�XQ���gϻT���?�JAg�%��u��l4H��E�3^,���-��@ծJ;�����,���R܉�Y�0� )���h<n��ŋD�P:ʠ�B��VމYw�E���pXPh'Z  �hX���C�7{�:�4"�D� X���w�I����I��^�J�������-�l�ߺu����DgO��w�ε�{��{)]��:��	1��`�"��&Ӹ����)@a>L
xuq,�P��}3�����L�aT�5�!�,���.����H��:׈̐&"�ﮓ:��tI���sml�81��=�=��y�ѥ �]XV>+�8�9r1�8XȌ�YV���׾p6��q�Oe���-�9��|D'���G>򑢲c�!˫�[A�+���H[Ԋ�%����E��FD<^�f���C�-`Ig�<^��M���nIu�<����\�?4��W�7����^�k.�nN�������B�e�$S�����%h۽1v�3X�����3 Z<��Lm}���3S�r��tҩ���`�d���U�d����@�.��䟌Օ�k>�o*��%�f����T2�jDs)�Y�M�x��������3ĩZW`�"�w�g
/� 3�Q�[�����E`cG~ӛ�T�0�������8�>�M�k�4���j.�>�s��\҃y������C�����u�ڡ�f�����Ͳ��C�{2wj'�QDAkG���W�K��Ѯ��;m�Μ���x�7�AU
�*Lt�9b���d�����ΰ (�h���  �3�|��nGt�(��1�Đ�b��,�D�n�.Ѽ��i�E�h�캚�!9FX��\���\��k���)�J�J)�ٯ<��3jf���������N;���#2US��A��A�8;3B��R��{�w��r���cN^�9�ݐ4CE�.X.4���_�Q
�@�w�K{��q_�s�>H��:s�r�>����oIZB'}���]�Z��8o�oj�mtP^����6gϟk�7w��u��n���X�q!WhQ�L�<�o��Ewjǈ��w��3%�8��f��	nXS^6������4mc��ն��K���ڜD����J��մ��E��T�Q�=��nl�p��U��1�Y��EW��w^�WcsQ,�����k�(��.�FZ��h	(Ζ,Ma\/j�0�9#E���]n���U)����0�n%Ys�*0���67�5����Q��.vd�?�wv'�`�[K��Ɖ�ϱQgF(�\�Ex2�B��PX�nD�N�L<Q���N���zO/z�	���qMuZ�bׂ�5�3��U�\�ḿ�lӌq)�$jS�@��*3~T!�y�ť��86
�T�6@`q=�-�s!y����F�i�{-{�qHZ~Ja�(�d\\d2�85A�a�^�v�<94�qmHm�y�}LܨX�;}<s]��vv���/e�;� �V;�KK��8��Op)�n�C��B2İ�ӻ��n_��t�Wl�ﾲ]OW}��h��zŚ��u�9yb\����얦��k���6�O����Y�r�2�,y��X�tR>�Ne�I�3M��5�)@Rșƪ�
bJ��bemUX�>�̉���&����'�Œ1�
)��M6A�]�KCyF���(o�;�S�)L�\8���9j�>1d�J���|�}��rGp�s��!�O�N?F��8�|��WM=���!&��7�����"�;�`�~��߅�-��Rk�2I|hW��N�-K5�щ���ک՝��lJ!��}u�l�b��=o�����iVڱ�z��f�?.a9n7�_h�����y�U�ze���kǵ%B͑���~��D
�Q��r3BU.��W�WK:�ꠅ��頼_M5�f��~��|�Y�����ɘ0�uT<�H8mԗ2�N��3����i����C�{�!f)D�Eϩ~f�L��-o{�ۚ�����X򥱻����L��@�E�<pw�)of?)�r;yy-#0܆`f?��8=���:��ej�fa��h$�
ND�vk�Ȥ�Y�&ΏI�(uo9��N�ܐ1���՝�W�v6�����W}�E��}L�;mek�-nX'U�K_�vƥ�餭���1�	��i����|3l�J�vONd�	��L[����)%ӊ:-��w�I�'[U�+��Y"0e�E�:Lތ���)��>�L�^tE�])�:�uĀ�a3hG�8�$`{��ҟ�fι!���󬝒�D���~5H�l,zj^�gTK���"&�s׵�Y��t��4��?5O���Y�n۴�-+eN^��n�������9������P<���7޸2��?bo�����G�b8��XN�Tk�V+�W��ca<)�Xl`-���L�� �T�e�E6[3������L�a�rɕ�Fl���TSiY|kR�	�ʐ5ⵄ⥎��t�9!y��+��LB��/��4e9~VJ#L��<��$�m�1m����?���~�2�NH���z}ۇ�i�S"���t��Z�,���0��d�q�K��~����9�1�_γ@�7��	�T_�.�M���y�c�C��o϶�̭O��x�Sox�g�n��G��[n{�`�oX��z��p��S �v��={g0*q#'Z����l6'N��
K:[���n���&		&�� ��E,��'g�&�B�(�(��oJ�0Y��qN��6[���ښ��7(٢.��3.)���:4���������^"�4}1$< ��A#���Fiy����B�*�3�7#���1P�1�����W_����d�l�u�!A�fO���:�Ut-�ʵ��_}�u��a(�Qɳ9ޔpg�:V�(hA/�:n�Ȋc�z�L��k��Z���湝ǯ�{�3������o?��t�����k[i�5+��IWK{�������q����x[txr�9��hΞۜ&R����|`�	�gr�s�A|�63�3@���|O��QM�U�Yq���t���`ڃ���q�v����Xe.�
$���}�R%�!ǖ�s\ja�3[����a��?�X�чSM�EC�|='ۚ��4w�	2"Pڥ=^���w��S�UѪ܍E��-}������ c(�ǟ�n�s��/#���ģ^q�"vX�E,�cBA���KKZ�K��^��8�4�L���7��S����{�I��g����n�����ǭ=�Qͭ�]��u�	+Ý+Vʆ�Â�K�{ㆮ��0��j�`�!���:�ew��1��wu��g�&���2�67�p<dc��Y���r�6+����</�-���٢{��D���y�g���R� ү�ў�����1���@�2ce�~A�6\ZO�Y%b�����{ɧ.�6X��s���cjU9?D�"�j�P+�gN���A$��G�8�wT~�\��Txjrr���>�*j��'{�������Qq�x/K8�joxf��;�y����x{ȁ���D7޸r��_����OY�����!��m����R-Z��C���v�J��F���V�����g>5a�a����0�^��WM�����R.7�j9����ľT�&��ZV�ʭnCi�K��3�A�@��0���,�d�/��,��Җ�,��)��Dڼ3\K�flo��B�q *�%���X�y^�6�ϐ*��M���وP�
CFBh�b7g�0��n��E�Ĝ܇ҕ��sσI�~ꧦ��9A�u&�9/2[�=�m����<ƉyTk
a��}'ьs�����rG��h6Z9vb��Ki� ��Qg8h6Z49��z��]�|ss��w>����^ks�
�}⎧������{�z����ںN�I4�8ך���Ѷg�}��hՉ�v�yc!Dm����)�Rq�\}3��>�^�Bȩ��(Ԋ56��`&���ht�Π���&`V��v>m��q- D��/�lE��_L�h��?j;fF)ty�DN^���A���O��6�'��6��ΩN���H�
��d�M�cY(E�)K����v$1�!\��S ɬQ�T�KH�����nsDQ{�0�uY�uu)`�&�v1�0&V6tN��c�X�O�*��Ѱ���ޠ���������i;u�
�a����gn���S�������7��?>���Z|ݟ~�/����/����x����+(K�&��+po�LG���]��v��y�7壘�D6�3�©�����Pb5k��P*�#/��mͲ���|�̧J)��ȳRHUJ�q��j;�1�-C�,C�	��6�@��E����h��{�Yז��ꈊzLs��̞T���3�*I�1Ρ���uf��c��9W�N����]�]���z׻�Ü���ٮ\�R����	�r�1��t�M�(�u��i�����4j������[]+[����Q;N����͗��h�;9>l��۞������������w����O5G@W��3'N����in��[7��E�v�>����:��~ �����}�mF�gt�T��.�<�Χ?��� TO:�dl(F]T�ļ٤k���0��&`��L~��ɉ�3&��E$'oz��=���p.��E�BB�f9&GL,�:*C�xT&��M��qн��on^��וJr�%���X2Ь?�׹�V���o"<#�����|Ԙ��Z�?�ݖ{���aoeg�26�kK�o�� ���ŃV�g�;E4���#���z�+v��!?�Ʒ�x���=D��k~�M������o���7����ۛW���ۓ@�X�܈�"vx������͸��|�T��F�ZO��R@�z�]�ݵ���|f	���11E�:���oR��!Q�IJ��	�|�/��5�����늶1�Y�1��yη�LEN�./Q�6����}���0��~N�0��-oi��ۿ�b��pNa��w��1�sc>!��(J�v:��6y���< ���
��;->?�vJ��x�L2ϲ1�p����J�P�w{p��w>{s{�����#����_{������������s��So�q�\󹫯��/Y��5w���[�~j�mQ{|����~��/���wƏiGU����Q��\1]���{�ʉb�if�V�J-"m�NLQ����N�����$���[Ln�M|���,^��j֤�oC�f	�㶩gy��\h�q��(�4 �%�[�N܃����#?�=���ȏ�HI�f_<l�V�s�K�dF�8�� �9����.��L��j���7鷝�س���6	�\�l�����R�E��e���(��IY�5��Xȭ�H���P���Z�w�k�޻}EsŽ�w�=����W���˝��w��_���w����o�f�8�~�n����qjcutzx���z���YW�u�3N�{���g�y�����~����vo��=��`���a��P� .	��������6ᬠ� -S�t�
+
ΐ��E�t��愫�&\n|(�y�Wz��&�	�S)��s쑊�&C!�4작���A@3��]��k�p.b���&RDș�,E;y�k����YD_�a��������[+��	�Bg�a:��o��X�|����Ú��,�T�ﶝ�{W#�Q����gvg=럍mV��b#C�#%Ĺ���-nV�H(\r@"6HH�K�,$�	�A � !���(��8��z�;?�U�{U�zjz{v����'��������W��{Մ�q��ѣ���EO��VU�*ݒ\<�[Q@X\۵+���0CceB�W�3$I��Fl�ɭ���R��^>*gO$���hddf�HrE�M.~�o��^�i[�Z�<���e�I����C�4;�,5�'���Q���PF���=�1.h�%�F������zh����XK"&t�@"/���m�_А��2�]Q}�MQGD�D���K/��E�W�ԡI���|$ȓ���(�>}:'�li	+l����Z#	�ॲ������Y,��PG�:]J��K�U�����}��j�zA�H��G����9�`�$�'P">t�P�lI��,(ݢ�IS�lH��Z�u%�S�oBu������ f=[ȹ�S�/|���$���ρ4�'��0f`�`R�TSHÅL�D�Jq����+6� A��D5����cB`�I�U+sY��(�y
ucB��\g�h$u� �WR��P?*�a�@�u��4;��9�� C$	3C��^;���`�Z%��P��,������/�B�Ӊ�}�a�t�~�!_��gb�'$�F3>DqUg��_��A�����&w|����'o"�$9�h�$LsT_Ɂ%D$�^z]�*��"��(Ġ��_v�����Q�#�:}#$e,[tLB{}�b��%�*IȾ�M������E�/LH��.\ )�����bJ2�?n&ѿ�8y<N�Z�
FNC[5-������a(u��E���8��x�ep�U_D�i(�Lڭh7Ƞ�3&l��ք�d�����R�cf�"�����+�2�5;���J���\]F�垅��sd��}�Z�_�����>Ń%�$�~�,|H���r#h#m�&�N��0�=�a��!,w;$5�ݭ6�+vOKܓZ�:$�:zx=P�g%�Ǘ�}&�!����Ɨ:'�Dj؝4���Ȉ$A$Q�u�e��qHڤ�݈o�l���y�}Q�j���^)�|1P�on���߈�I�e�쓳��`t����Ե���$,���|���b���Z��w[O@��Z�yh�PYG�*k5qKP՜%7�&�/�<=l$L f�����%�Ђ���V��q�q�Pd��R�}x��5/H�x��$2�8k��*'����q�U�4v��đ�L7�V$0r��-$�����m�{�( �M5�����L
 M��TK����#�@�
LIe&h�բ(1^�ܶ����F`5;ٮw���}�Ң]�o��ە�k�B���ۤmc�7�� A��oޯG�_~~�?��'�~�����I��\��]�>Eg�S����Aq�A6��<B�R�����?�䓿y��W�R�UIU���O>��w~�R9�Jh4��.JH�>[�\A2t��Z����1�u�"�J�
͜K4��ƨ{�&p��S��њ{i�Φ�i�X��y��u�S6��T��>�|n���k��Xa������_-5��
�@�;���{(�=��r�F+�(6�.L��t|��͕�F�ïK(�I̋1���l��� ᓄOt�ٞn&zIz��z�[��F���|�z��I�4"�dgMs���o=����:���b<~c���v�>�0/���]��X�F��z��'2�2�vY�ב�2�% �,y��ƥ��:�.��y��2��WweŘ����M�Zv~�4e�KR�pz�!cf�f#0���s$L�������Ҷ���TM�r��)aI9S���U��(�߉9�7�@��E+�L���O�E��v��(kk������ҍ^D�Ϟ��Mb��r��e:ύ�|W�2K�A���H��<�*�&���bؿ
D�H��x�g���$���^�9�ƛ���H;m�MYzTe|�F(����d̝����a�bFf���ˉ¦҉��L��W"����N�)Cʖ�P�v)뤬���|�����+��|��׼������n�%�N���&Ν�;/B��N�|?љ�T��0c�����D����̩+� ����H��fLnI��&�Z�� (кo2� a����:�A������,�{���ܢ�����?>��S����떂}�������?|��Q�[z>N���1�b{�*5�!s2��*"R)j�'��b�~��v�Lc]���c���-�9q��'evQ;�w�~��V�LsI��/�'�hێ:��V �$cn:͊v_IG�<���V��� ww��(k$�A����3�aK������0Q�D7C=�τw���|��=�Û	mgV�/H)�LLL�=r��/���9v��ۈ�Bv�ң��S"b��hvi~�j�>[��x��1Wh"2C^��mA��r�1j�ʎs;�k�QG�H�K���F#�褶p�ɮ8�J^H֙�S�Ga��J������LKnE�|�2f�%�F$(�k;�e�ۦ��u��J��󗤺��-��k��i�Ӽ��n,ȵ�����p��E(�k�����b���;�Y�!`#��>�j v��|8ۯ��Q&�o$��h�Qy�x+"7ȹ���Q�V�-�7���ܾ}��<v��^x�O6���[�OO+��'��F-�}�+s_�K��h7�<"d<�2U�*�@sM7\(�y%�:�� �I��u��I�ܑq���KA�+!gn�������a�0k܆�]L�2W�Z/��Z9�K[F�Y� ʮGm��	[� 8|]e��i:�U}�ݟ��M���r���3�C|��Q�r�5�g:�	�`^DѲ��(��qeTF��
ɭ����$���x��M�<@�ve���o�t	ig�.�Yv����B�le/珅�k{֑Վ�g^q�U,4���E�:W\_��5�z��}tٟ�A��Y�.��o��Q���j�\~�#���FGG[��M��?}�����O�����_߿�={���=�3]x�[7��g�V}��lt����X��iV������{Դԉ�d�ⱝòt����p�t�)T1PqUe��E.�a�P�]>�9]h��k�/����IRvS�	\�)��C	Fl4��}���FSm��n�.5,����r v��͐�� �1-@�7����/
	�Ur%��@q���r!��mvg�င���+���(p\d�G"�*V<�Q4�rҍ8m����92r�Y9��t<����y�N�8�nvS;�l]�#|����,;?x�F�V�یu�a�y���=����x	ҫ�j��c�=V�8r !G%�T$�2���E\D:DR�}^�х��l��,�����7H�������;S>*��r�A�%��|W�D����D��D�8�@����^x�"�v�DĘW�	Mb@�}�����d���Í�{n�̙3l��>�R���f�:���7>UK㥆N�D'�v3*V:IAք&E��ɉ�<�D�I�0�x9j�Q��	���$uǪ�y�J����ߝ9>=���٩)�N�T��s��_a��W���T~�����ۋ���v��N��u��g�u���Y�_��SǻuuvV�LN�=V�KH��5���|���LMIv�<:=][����L��Z;Sz)br9fzeX�>���
i�d/٘�Sc�gV�G��2�>g�k$�s�ߥ\Xے�8M!���Gؿh;� a?�}��ӄNT���+�J�b8�D������_����x��x��ָ�����C�ML�����Ǒ,�-c��Eh7@�}�СCOMM̓���AE��y7HV��z��M
RfN��Q�^�a���9�_fl�������M�k6��l�������~���͙����by�w�N�=i٨2]��S�ɖ��,�-���I��2�!&3���]#��X�ZjT�� ���Qm��e5��"������A�w�n���V�&z?������20��(����k�g��Z���R%�@����Oq�ʝ8��@r���
�U����0^,I_(��r6 �
��Iv�����;w�Lϟ?��8q������4<��U���v�h6Z���.^�����{wף�0ȵ�H�E%��@0�SβD#Y%ZF�8 	��L'@2F���r�w�Q���Z����DfQǑ�*"IϦ�OQT�<C:��O
�Y����R)k'i�J�T"ɡd�h4�������������{�l	oA=s����W���.�-����إ��y%޶��l~����6ν��<y�d>�1	�t�Az�F �-�	V?�kl�0ξue���NS���N׽�� �7`+ ���V��V�]�q������e�!k ����v��Į�I�ㅙ[���/�����!��������GD��F���w���p0�UL��:�;I���ή
׶/r�'��ga�dgaa�llafbbj�p8�R��hN��҄��


	*2.,B|J�?���m�X0g�?x����sJh PK   �yDY��� 1� /   images/1e4fa634-4e77-4d97-9022-ac13a26749b2.png�{WS[�n=�(գ�Nh60B@D@�J�� `�����&)��b�C"-�sw������w��1P{�5�,�|�����jk;�u�ܾyb-�ؓ~b?�����:��!�����?��î��<@ �Z�7S��}=��g=o=��s��?r���pq;g�G���.�h�t�y�w�� ".a�J�G�V��oB��ϝ;����e���ֺƽ��L�"����ܩ�H#;ҀS�~�|����[������>_ر�t['",��R�WF�o��r.�mo�}�_F�X��u76f��K�A��� �#�}���ٿ�4���Oj�K�u������g�]�ߥ�]�ߥ�]�ߥ�]���ҕ�`P�a���Vna�����Ha�uvRا����nBsH��|�!4���?K��Y*���fٻ��C̷�C��R&*7W`��i_��_�ή��'�0�^�D�O>���@��hx��UzDh���ܖx{�JD�:$�;�CN�l�ՠ@}X�n�����=�e�ՠ#����O��E����e0"���!�=��pW-I�G��g���jǤ'��"y���B���x����\��U�$�Q�(@��&�n�M�;B���!���3��P"l���ƫ!a��c.�d�p���g+�ө�2L�@��z�~G�r��{+��;��3���ʥ��Ȥ��/^�	H,��3�릍��@B�ukii��|���Jo��j-=�+�G"�	߱:���F.�z�b��2��?5���$��)C�E4�I�Ͳ�O���s@M�<G?�i���T�p�X33� ".�}N�UE�YCv���W���x6\;ŏP~ �÷���J����RNX�`sg��Şr��@f8ܬ����*t�hX�l�˖I_x�g�T�'S+����v>��4�!q�c�L�V���-�!����~��)�o�fm|c_��S�~aD���"�Pa�Ls��.� ����l���?��L~�}�=au�OT܁�W&�p]���v���iᲿ��x9z�6�ɸD��d�箳�*�~݁)��J��Be2����ȸ�ĳV�a#�,r.�_ic���{��J��:�/Ļ�έ���S~�]��7\���ϒ��Q�n�����m������2V�9v�6~c�AXkx�]��;r
ͤ�_Ǽ2� �r0iX{�(f<��,s��{Pna����ϯVF��7\{��[�!��K��k�&��1H迼Yy�O���
�����N�h�eQ��5b�9�)������ٛb���t��le��-ҵ�)�?Fsl�z� n�^OYx)�)�ț?�i�-�K+|�g�c�Iځj3@���*f|��yg�J3Ʈ���
h�Įqbe$�,�{�P�H�P�)��at���2��t�.+`�Κ% ���*��FF�Y������ǁ�q�ɗ.*�
�KO(|~)Pv���ϾD������Fd$/���[���U������8�js� t��gj$�	��]��ת+�±�����Ovlgv�	�:&'���0������W1d�܄�ɡ��tۭw�F�/|l���#Fn ��@!wu�G�8[C��6�H�Q~Å�8�Ϟ�J�Z���c�uY�\�}�eLdл[�SR󪁽����+����W.�o����[�5v�{���0ͫ�	bd�s)
��,�3f�Ӥ 7�r�_�z��ԅXy�����owva�%e�0:Sߥ8$-�=6��Yj���?as-�^�J����~��}�d��P���^�U�(O>�Ȉ�C1�]��A/=!�I����!�o��F:�����[���|8A�_		�)��;{t}��j�XR�k����W�|���U�Rc~$�|n`"�=�'�Ћ�������v�r��-�f�?ߨ�R:B���o�Ȯ!�m
y��^�U����ƕd�U�9OŘ�+���n`=��$U8U���רR�ok��wi�����HRx�UE���5��R�:��6���d��Ʉ2�]Vc�tuv�x�zJ���vu]�p��1� 0�S�B�Mo����ȰX�7_�; ��hy|��~����U���~T�W3�OSE���C��I�C~�E55j�0�Q�̚�'��f��Zzzz�q0�5�+uvgǲcw�4���MT�U˷K�M�^G��}G��ն�W��(�+�"O)��v���j�H��w��ʸ�O�0=���z��
� �{W�8���#@P�Vµ�V��J5�S��tZ
E��ڹ]�:���P��e�����ɴI_�K�%^��u�6�f��\������� "��������-��i.[�3�۷ⓑ�y�?z���|���� c��w�(	y��@fBS7ͪ�h��v�;e�L�+��}�d<rȷ�+�7�xÀ���-�kh��s/�>��Q��A�Ļl{$�5C#��y���:!����5��G��f���Ak�x4o�7wVߨ�7x�ʮ�1S��īu(lK ���X>�Ҳ�h�/\V;J�S�"��I1��I����G{�ݯt8�q��ۂ	2�IO�v�D���k�!a=Z~�5�Vu}-��#�~y����,Iˇph̑J�����L�G?�]��R=ގOw���Y��]77 ��0(����z"��-i"����F;�S}��c�*8ޥ�V)1�Us3x�Aw�9*�|XO�"�����dA��n��(´z��O�B��v��x��^_)�)�(�?����`�e����"E�9}�{��-N]J�*-#�l_�{ߝ�ps�a9=�2�#V�Rk�ۥ,�>����VE\�无jV=z�Z2����컫
] �s��w�@ڡ��<�|p�uj፟�J���o���|}r8���SW��K�_�Ɩ���@*����=�����( ������T�R�m$]|D��ήP��R��T*���Z3*q��g��G~�Wm�,ٖYd��C|q�%G�*{g�vUQ�y�}�W~MT4 -EEˈ\��qN��- �/�[�b�ȟ���eN�  |_O�� �	���<�" �Z��g�jh���1���j�l^-/!�(������`��?s���D��uhG�3�2����#;�������Z���I1��59p�����E�y�+��.�Z��D�'l����m����Vn0b*\ʮ
b��}�EK��T�-wi�0�
0f?y���K�1�ց���Q6ͫ����z	O��P/��͌�����7�(�>�y��ح�Z����(�ֽ����&��±ց���4��=_t`��!�M�wn�ᬉm�Ea��DMC�U��q�b�m!��ѫ����>��뚓S�S�mšf�e���y�!Lk�G��}�;�:�ߋ5���̎����~7�xSc��-i�f��ä����j����������e�pU51|U����4��� �H�6ȃ-LB����Q	W�>�o����j�6L���m�x.�ʙ�%�`0������+/�6�s�*���/a��$���֣`�N
>���)c�O�<6C�8�+�c��|��#��?ײ1���7��y�M����uɧ:�����^�*�8��Vh_D��5�N�1�����:����6�+�YNU��qg#X�Cݻل#I`kp,&��9���V6�&��m!�����|U+%�47��WOO��}�b\O���kIu��%x�S�е޻��'f�.o1���
��B�w�,H��}�����۝��;δ���s���:f�}�e�������`{�w�����+|}�C���;�M�i> 
46\? <6��\s�]E���p�����N����mҏ�E�w��l�|
k������+�]҂��-�Sc�^�1S�{~38ׂ�*[a�*�ܜ�a���������W�-XꚟǴA`�Jp4F���$���r l={��^�"~����ĿP-��i*~�1*<��`�˹M�P� `�~�O���w�4 ��R*���'R��V@�5�i;��c�:^Ե�p��Ք�!"���`?:�ADؔi�
��Iֺ���UYchLZ�f�Od��M!<�~� ߪ�n�~��&i2�����j�!M�
o.��ƹ���6���8�NZ���n���a
�y���=�(�6��zu䀐�#���皴T��C�]=�IS�Z{�����q��$N��fs���ҩ(��L%�3����04B�u������h�"���~�!����;�\������?����uUY�d���l��x~g:�6�D���׮��������s�_�x���:�?F�ɱ��3t*�4��ݯW���Y�L�-j%�?U�C�%�ә����*���I�	K0�-fsZ���Cy �J�?2��[ K�:uu����l}ctC���m8)m ķWF.>}.��B�.�((��ݹ�2��{	o����W^�6x|x_Q$o�4g�b�T㱳Q'�5N��?����+�'R�Cσ��h��X�˩w{�'�VME���NUOQD�șz:8C�:ݠ���Z����^�$&2 �ֻf1�����>6�щ1pqSK�:O���?K�ߨ7c�Y͵jY$qb�w/���G��n3��Y�/?)u?��m��>e�ӛ���Q��8�Їa� H�`'`k��"���Ԡ�Â���ţ�Gbd�_�l��bl�٢)f���սAIR�1�h�e����/c�.=���L���7�$Ɲ�v�̴�*�w�6!|Ɵ�Z�#%�+���pE�Q�wQ��WG�'�	�G���H���n��>OM@j_�; ���b���޶ �f�C�2�7�:��G^^��ƀbU�����uuZ�"��c�8���-�=;)Nʾs���^��C�~#;���}H�N$�z���Y��V���-P;����<l9��Y1
�&?@N�sY���!y��Eʙ̩ޔԩ�,/}��������rV�I�@2�s�e,����S����ɽ�|������=�俾`��L�Z7u��&ҡ��RT-�w3t��7)q7
�Ĺ�L��>J��N*JNIu��x��ȉ"J��2�[dX�c
;�D��<N����޾�'����+,a6�Ҕ�� ����|���'���`�E�������5'(���>~5���j�^�M�m��m��v�fy~���.+b		���Fb>�����G/�-���ut ���h<���skW�<6}�P���D�����@~�M1c�����K�O �����w$^�c�M:5�3f��m�%j���9�vpD/�_7�I�����k���_�`T��E�R��'�>`K%LK>�a����7���3��{����=e��nI�;��iᲬ��"sM#�R*2���D2)8f׷�t��ے��=l�кkm�����zaν�zB���W͐�V���]S��>J�P{v�	8e�xD�W���\L�11(i�R{%�^�z$��a���	�5w���j=�!˪���f��¥�� �w��r���kt�'�Hy�-�`e��M!�?
<y�F_(�1o��}F&�uo�W�5(ɻ���jl���\6��߷���� \��� Y]���b,��w��S݄(�tAI)�@�rz v/7��#2�8!*҄]���@d_���7������1���y��o�4ړ���¡=X�4�y� |�a�Λ$��%�E^��1�h����W
qn���1_��y�\B�tФQ�1�S��&"3yw���P�(�����瀘~�k�T2��3}
�%�X�yn0��m8�T�� ֺQ�ۻ�;�n�\!�4��yp�<���ާ�i����hW��m������kf|, SU����°��*�o�;�� ��tEn3A�����Ġ���pO�ĵ������ZME�������F�@);o�r|�,A�ה��;P�gC�u�	O�ע��m�����W�v�"xOԔ9R|�j����#�ܜ�3�m�E<QJVf��䴺MP�YmP��26���=\��g";r�&[s��y^�c ��ν��[OB���7�oO����0g�����;� D}پ���H]1�3x뱘���2N�[737]z|�����kV� �� �yx����Ԟ>���9�8^����bYv�<����d�-�X�nR"&�rk�(�1c�rkfF��z��0���VUE�u8�����q���2g�⛴;t(�h�<�gI�?�XA�X�5��z݃���!�w��	4O_KYN�ٶ�t�V�͜�W}Bx2��`�����8�05<z�&�}��o���x��<az@M_��''�CX�ލF�D����ˡ�6 ���1�y��,����<0	x�� ���~�n��	$�F��ST���M�䖒!�-��ێ	>3e�)w݀�� 4^Fْ
�k���#D����R��+���g�Cx�p��w̆t B�>HX�������ޙz��,�H��jpq�I^&�M���Q�{M:Jg��l`,�Փx�f�j��Z�&:.�_]x03k�ؔ����>� �l�;�r���4���^I���S�G��]ء�W(C(��~�+�V�p��'sq9E��R�]f��`�)��l��,�;a�21��U5	P��p��BE�X�vkXG�[e�j#� ���aW�UCI�q�lW�(�;U���������1��K;c�I\-eI��h����߯�Q�P�=Z�IK]o�ʸv�1���p=u�6��"o�	UN$~e�v�	R�.>�ї��AV�\ t�J�b�go�BC����cEws�0��bj�l1^��7_m��ޡ}|.���KgL<:c,JGX_:�X8�����%����!ǳ�*\��P�p���jZ����Z K���%l��-�۾�ը����Y1܎*�݃If��-��'~�vXM$�
�cý�+�ﷅ�-`GE��N�F���_�"��|`}f[5�y@_�J��"�DUs%�����2�X}�J�Og�d�H��qs�H?!�qH�ִ�b'­�m���mB�����������gx���}�U�1n�v�3��qtʖ������\�ݝukѨ��tj[�ˎ��&�f��~�w�Tr�L��)@}�K D5ڣ�˳]�w�j��9P>m�W5�g����&U>����%���+�5{��wyβ�
l]���k��)sk�n�`ݵ��WQ�<���Vη��m��6�(o�iU�v������s��w7�:�	�S�tw��
HP��[�3YS�
r;��@���4��Vp�7��%>�]㚣k�ߝ%, q���y��"�K�4�\u�C��� H1�`�BM�pOb�VG�8=��j|*.�p�\_�W�nķ��rp��(  U?��J��6o}.��I{pv�;[0gZSF�Z����xn�Q��ٯx�M��?���k 1�hr��Q�#N��J�k�憪H���B���VΩ/o�ۖ�[[C�q�/�"�ϩ&qc�_� D�D7���W�Y��5�N�D7�)�e\��.&K�(~9hݔ����g��'� Z��^���˜CqȢ��Ҭ��rV�B��W��2��L;��{NސP��H��_��-)e�d����iX�i��!�S��t�o���Mx������G%* �#?�We�Y��r�?q��L��v�?$
V�GL�㱆C�mQ#�$��8��f����ͻ�z����"�6���|@l�q��~VKG��FR�)� 5��N��X�G��=��-�l讳a�:�.�9�_�-�<��+��ZBE���E��,�������h���p�d�� ���j�l�@8�ﺦo;C�Xe~<�d���G�Y�PI@|�C����|?�2��\���`d@�13�Pƈ�nR�������>�t�Y*)��<������,��m�]8݂�?l1_���Me����,�i��m��T�d����EĳS��|6|	*���y���j�wLe�+=u�G�^Ñ,}�b�C?�e8��Y}�����#1��9��%T>���t �g�$��ܫ��a�B�z�m��a�C�c�m�.�0}dg)�Į!d�������Dy���SJ�:/��Z�eb��U�/�1�.�G��%G�z��r�G[���3� �T/^6*���:�~=t��[�s�!:��7��I��u�W^׵�,*�簌��.a<�*q�RȬo6���-��`�I�UbR ɻ'����Yf���pByJ'B���f�r�C��_���O�����Z�Z�	_��^A� �۵���L�� �^�ZP5��
Vj��Θ����%?���� x��Bf�jRqqq'�1���j<�N�n�~�Z��(����� �G֩��N�zP\�s91Gs�hA�6zr��t%�/���k]7 9⪛�r�*Xe�IT�I��.q�ν[U�3K���䧹6\=���]�v����*1��&�O+�e*49��&K͘�����m���	�{c�w/[OOxzZ6?3�R�������П�̼�H4&�/Qf3_�Ld���vK���ʿ����I���plO�N�)�N2fw��B
x�< Z�����0P4��u�Y@������ʓ:c4=nYq�Sh�~X幔���BKHZh�9lo�%2YH��P���~R�m���87:ܛ�p��g
/q����!Q1�b&n�{=��|�2WCl���\���ߨ��,n9O�ho�݁)�������gv��	PG�_*L�y�'��wy
{*��'�d���2Y��~>ٚ�0?-fr�{%����l:�6�L;U��qS\����E�ɫ�����ˇI�M��f��"�Ӥ'��F�0�+D��S�O���%ƑE�����+�.k�r�� -w���_�(�w��4E�߂od��o;c8 vXI�:�j�kӁ6���s���mUѢ6������S��W�������}F��g���}������>�q#��N��KÂ
t���Պ��5/]\T�&�q�(�n��NP@[cJvo.[��`������^���?���h�4��f�E��dv3@��N�>�=���WJf��j[g���=_���7��#��2����2� ãqa	��րJ��-
����6�ܤ0@V.�M�Y۝DxX����d���j>k9�����C��"&ؓ��D����[雛0�����Ҹȋ��\w������A^>:lR�W��Ћ�ֶ���w �Z}܇��}M�#ږQ�e�#:l�;d���r�
��mJ�צ��W�!~�:8�$|G{�=;�$�Uŋ��q�W��Ek�;Yv�LŌ��;�W��Z��3��p�Is}CpM'U���o�V�g�(m���S�ѕ��}�N�����ap$��J��`�R�W�������B��3'~>�ʽ$��>3hS���Ee��6U�}�%�3#�aҪ�v�ۮ���t;<�>7���Gx�I3���ԡh���vV��___W��~g'%.�=�*�OS��"��O^z+�T�����$�R2��o�m�����qT��~D|�*���\�� �&6y!��V��l�@ZU���@�R.r)u�➯g�ջ���{��\>{�`���'m抲����g�s��KQ���=��+J��t26�B#<F��~���$u�Z��M,�ш��w���ڱ/_�btb�jd(&��R=������-=�����~�0%�q%]�Gd�!!�aҙT��f�2�Ď:15��E�8�2���jjs�+i�8�R��5�Y�!B��\��ORm�D]��t�|��\0��z��0��%ð���A�+���TKΐ����ɡ���+���@��z������~��$�Q2�s�j�H,2?�r�Bypg4�eUc����9_3��$fR�����g[�B�s.=�4=��'��h�>���8>�8vh�)����̻���Y������ a���������+ߦ5VЫ5�u~9:.���|L�?|=�a�c�s|<O�ұK��#�d+�m�
�_j�oqc�h��&��p���3�^C�GA![�w��l�b�7�S?��zl1.�w�,�Yuh�9v���ވt���F���m���K:�լs��Df����SJ��q��0�P<::*�< �kQC�9��5r��˥)(� �[�iP�B�XǌF�����\\�]lUO���ff#���0qj�b��3����%U�I��$�;w��|�F��ա�K������_��OI��	i[�lpB��͓n5u/�W[�|��U5�LeydN�~�x��S-BpV��tF�Tc�ݣR��=�t|"��E��Q���4��\�"�@���R�R��R���G��}y�~�{����E���\����&A}y�� s�#_���zoNZ���ؒ6�We��G?�z��p�Čq�k�0!�
�Ϸ����Eb�Ɍ���vO��xr�Q~V��۾zA}kN-E �z9�I�<U�05v�u�aX�Y:֢5�ҞT�����������\Y� �Pz��޿�����-9����5�(ώ�"���~�Fz�{�;"!J<ȡO�/α��+�ߐ���~���YD=t6A�;��v_�8�:/��/$.�����#���J��"ݟTd���T��M("�3�7w"�a9�� �  �y��y8dcv9 �-H��gU�&�a�*J?��<S_s9Tڝ�<D(n��b
��-�[-J�v}��m?*6x]��Y��M/~�O�ek�SlT���/h�,��$-4��$��
�݉��cV�5��Q_��`�Ev��|(+��K��M��T{<�|�;��=��݇�A?���eDc� �LB�;�<W&X"�/@���=�'�9E��Y�Vg%lBo#�t�Ҡ)��H�:�I�\�)��s#��tǈ!�*p7T�Uc�������ä�U�M-z{z���2%]��<��Oޔ���A:l�q�G�@ɏןNu?���''R_�Ӡ���U�I(Kl��*���rD!ͯao�~"�!^ �җ<�q�\bI���h�����(ڈZ��X?�F���Y�$v���Uq?��:|�<x?L�jն��0Vք�����J��Abҵ�Z>��s����p_�0�����L��2>�j��'�0�%�@��!j��v��b��|���t.M���C���?��e�R��X�⅟�fF��!_�_嫒s����#8d�&�o�7��?��WF
J�v��<��]j��VhjB�#�L}

:�7OT�;u�%P���ऍ�s|���{�e ՠ���Nᶄ���h}:Z��s����U�*D���Y7��\����2�f�}1^�d���?�k�>��U�X�g�p�'(:V��خ�ȴ�o��}5����Z��֍z�w���B�r�ϣ�u}� �6i��r8Ϟ����D������_^n��((���!}�ų7�#�5��m�P\l�x�m}M�k[��:@����1�H��]G�/�ޮ�_zJ���1ƮcPcF�1�Ӿ͒f,vj�|g��ְa:�<�>>��<��ҽ�ą�0,� $Ʈ�Q�C!��ݰB��*r�pn�1��7j�H�dA0r���0TξO�țKk��:tcl63ZQ�L,�����F�T�i�U	���8�k�� BЍ�Xk�3z��E�Ͳ�F�ܮE�Mb��\��P¶�r͖����e(7�PE�PO��NWm�}s���i�p�Oiӯet����Ep����az�!3��j"�&� �Vx'g��I��uH�-�R�7����9��#9��ӗ,���z���\~_�]�\�H�~}�ml�s��^�Ż�^���\�H��@>g� N鉇�3���P�9TU�W�*�&��_D�Kg�M��y�����N�
�U'�9E-�j��udT��>E3�1ZǱz4Ѱ��	nDƦ�,�2Y�`�����vҲZ5qH�
Z��kx���ʩ�*���CSRN����b}�Ěk��.^�U���K���u@.oJM�f:��aa���������:2�f�kn�wA#$z��+K��?�.��(���OƋmǾ�����Z�=�k8�Q���/d��I��X��� P&K�s;׾�U
ށhI��4�u�=�t���eg~����({zVf��#���˭���.�« �g1u�[��%F���cXN^�~���4F�[A��-�a�pȺ��}О'����IYyQ��ϟ_@��魰�#;D<z�a�lg���.L��O�J�^\���� �򳚾6l Q��:���|��2�)Ƥ���r����2TH��sţ�O=X�b�(�D�ܝ�8�I�0�拑�tҕ�`��_�N�<����[�P΁@�2C'E/���.�K� �'�p$����îH<�r�Q�ܗd��7��D��Y�y��d�)V�U��g��u�2LI���<�r\�||�U��j�t��%��qsz�--��~/��ؼ�P�-'�޿,1.��I�ނ+��:�e���^�l-$N��B�o�o�����y��MY������|�A�\WG��c��f��\DW����H����6b�R��>�sS��kӄ� ���o�O/�Y���)��/�;����J�ϴc!�e�KX���IO�!�6䯮$F:M���6b�����ڦ�y�bٗ}Q%�oN��S�@I�`�LȔUl�����Mnt��iP�[�Y�bϖ��Q�
�U�z��ö9��T-Kj,�5t�zcw�i?8�
���g�]�����&�
\B���$e�dK���%ØU�U�*�e�d���6D��jX�:$�J����3v�����c��/:��*K~�Շ��Q`�
�������j؛�7P�Gc��@	���A��.�I��}7��䐰D>�	�	w���sEUSVKXă�*�Ϙ��vp7��bSŤ��2� 
�U�?��pps;��@80�r�/����o
?0�<��"��]���p���T��h�����4���۟��o��eOlF���O����oo�t��ɝ3�����3)�ʎDp�C�w,Z����	�k�|�2��'���N*;G�n�Ь&×6��pecS������f2m�V*=�'\:�d�?�o���'h5��Į~3v����W�D�*��Sw��|�����;*�xo#�-6j��y�[�����_%Ө�3[�,�$��e�T�i�������jv-4��6��Z�CA��!F�`�L�sUa�:k�7����� �G]��!��Ấl�4���j�-�,�� ���(�;�Q�q$=����1���a��>�8�J�����ܫJ� 
\�<=0 �U]EO��P�\.�w�5�M�s����N�p�3Z�m���m�-/��ui@џ�D���7Y�����7睔Jt�7���� �:�ɑp����D���*����z��i��Gc� �w�����aT��ZaP����n�=;�����l�/+3SҁI�j�*��*m�.����{@�r�Ο	�Bo�p��<�r��F�*��&��8t�o��o7\�~���|StR)0��	�qPqc���P�&���@�kB�L\�d�A����ʽ��ɵ-��l;= �^���Sb���O?�Y@����G���;�M^)�F��-�!�93�f¶�pZfn ^�+YK6�͙��)qbT
�����@�� ��&+��1=Le�tK�c��`�a8�t�qF��j�t;����)}fSo2Q��M�i�v!���h������ivh��Xv����$ ��á>���@%�{Eo��|E����ްI���.c�ش���ii�-F�'>�sO7��ΐ��;����W� 4����k������b��G��ح�ʱ���e���2S����h�e���T�c��?	���2N�ʀ����E?b0�ӿ2�#���p}]ʦ��9�!Ʀj���yϱ��hY�Gwi�V�"��W����ݻyLr�
��1��� !�Z��y�5$�/kA�O}8�þK��U�h�{�"O��\�^��@��/�v���YF+�W��-��@�|O���o�0�)W��?���D/7��|�)$VP�Q�NR���Tq�-�@����`4�ی�3��(���������U��;�F�C��)5�e��a���\��_��8���иӛ�meUS��H�貓����)f�`�TWNT$�o�I���l� 'i?;n\H�o.�s������,Z�W�(4�8��|�������8�F��h��svY�xe���r{=n:x�m ��ǰ�3f����H{�G� �D��p�~Ssi��U�����l��p\���Gq
/�V�{�$r @�i��^�:@{� �^.�zC�y�2d	�����!�����n���+2�ƨ�f,�� ͨ��Lf� ���t�cuUG8߬���응|8���B��e��-�7���Xkkc+�p~]�d�@���C�I�lZ��	�m:Hc�z�q�'X����s#ݧ��������/[�tg��!M� a�W��7Tw}}��`YF�n�m\�@��sٮ�#������.(Vi���]q"˭��jO;o�oy���J��l�����1\�K��'Ϧ����˄�y/����տ�i}I��8�cO{�$�J�B�D��*82܎X1�C��u�G(�a�X) ����J	�3�{s���5
�S14 L��h����/V5f;��1�ڊ� ZC
�%r��0=3�A�*K"��m��$?$��o�Ё@Y?+"��%���c��S�8��>�K�t=J��gw�����	Iҗ����&�n�ͧ��a ���^�����F.�L>-�%�XZ� V��_���:{:�o,١�S�>r��w���9�n��zz��q����ūs�g�:^5֪��b?~܆D ?	�H����2�j�"�đ{Rh��,Q��'��p�f+�,��>���M�^<n �B�F�h&�Ġz�ꯪC�8������M���2����i�(7��xO���ݖ��v���o���r��:�ϟ�6�#K_ ��Ndɼ�����u������ܿ�K6ɢ�1c�Q�[|���[RWW����K.�+�݁«֬�����}\�)�S'��r��cJ�����r���"m��>�֩l<�So@Ƈ��F�1L{iT,���A��WΒ�D�>�贕��ěcm�c�m����L|-�t�+m+�(�7!1m�Nd�J�1424�I7�&);U_�U^������m��:���5@���"�|S`�+�����dAb/x��ɻ�d�\:v�w�%s�Nw���}
Z_NS�&�8���<;����h�>�<u�+��9�=�r6U�����L���Etu��-�"�@�:���ʧR�0V�p��c��#�m�Z�DҸB�a��ۙ���"�9<Ȕ���@��#��mgxқ�@���0R��B�J�6f���{ �қ���u�]��Ɔ}D���N̼�Y�T��5b�_i�XH.:�{�,�]����S�x��odk�sRgt�BCC��r�VD%ߵ��q����x��A% ����̼�{�}�.C�U�4E�#�����_Y @je�{�8�@���Scl��#�3�/�N�~�{���X�(F��8z��(����f��ڷ�3��w
	JaE�U��5C@l?JҦ;�B�Ї7��([H94>�����ȃ/2����`hs4C���~o���=�k���=���`ɧ{�����HFh����K�c��z�-�:��	�k�����$*ѐUiO�Q����Z�h%���$;^�B(�m�mԴƛ��3���Ȩ�-�	�Qt���7��(�vY�gQI���K�O�H�Ѥ� �	�)�ֹ���=!7"ҪJ$�V���ceݜ�_7���
c��r���;"��$�B�9�M���#���(Q�a�7���c�Q�&Y[�j��>TR7&]�v]v]�"�$�9�������O��}�ȊD�{Pg���3R*�7���-���9�ߵ��j2n<%ڑ]T~OC��=��-�-��D�D:�2���=�olp
cS�1��oS�����Q����j��h΂q`,~^���;�F�8���`��wl.f)L��28���;���H���d�x�p4�CՓj�g�8Xl��^kjH�5[l&����ȱ���Ծ\t"�\W79'�2^$}h�U��!?�C�}UP|G��H�NH�]��� ��m���9���/[���5=_����q�ɹ�Sl�b����>//��ə��+��nL��7���7%�~V:�8y��'(RA��`��ZtV�3�c�*wk4��J~ku����,���p�Fo/�l��x��P�x�g�r�;`P�̮�o�$f���O���dX؇>ۜY���hF����m��rc�����#m0����K[-)��ֹ�B�������.)z��Y�=g�㷨چƶ�>�b�Vq�Xd�"i�-+**Z�X�ax����(dI^y���[[�]�k�g�N���f�lrN�w�f&U�Ы��bT��ކ%+�Ц���Cֿ�ʓ%�K���4����ܚ%KHbLy#ƌD�;�F_Rs`<���BL6�i��9*
০��K~N���>���,�Y~ɶ��<tp �#�2���.I�VR�����<������@�c���s�g�a��<~c����9��H��BK1��s)�G��k����� �t����<�!��\o����Ek�A�^�t�Ԟk�^�sU5/8��Q`;�=���-�r��O/�N����\�͙X�)>�1�˪�7�zaDͻ�_�5��e���F�*�8��X�V)#��}>�<Q�����'��Ri������N��@I�W�=aL�����{2����=l)͐WV�x����4c�U�q�����Q���E���^�����{���p;�[����VA&���b��!RM�d�����}p���`ڡ�3���qd�/��1L��|�7*z�y*�5G�R��^E��:i���s�j��E(=1}ş&Қf�z�/�6�_��U���1��U���W�W���HX0����a>�Nsy��B�C˂W�2N\��7�-�7�yShV2���&F��)�S���}���p�D�U{�fbَ�@ :4��.�zX�B"}S߮ �b��FX�1����s{1�Z���R7X��#Wz�txT��hY.ed�&+�NLLL����57:6�(�J�� �4w������UykS�a�Q��n\_ΦW��3O4#4����ӽ����%�S@�����>u�?T��.��ܠ^�Jآ��� ��s����3������Θ}��
x{�'{u rJ-G/3CK9��Hp���������-�Ve�TɾkAY�6���ȖaP)w	%[�d�1�lc�(�#��3��9�]���~�繾�u��:s�{;���u>�|��U��i���ۜM5��K��zJ���4[,t%�PD�U�J���CvS��|��{��k��+��G��Wn9��Z�j�h}85,G}\i|G!*?�6Ｆ�aH�|媉a�Q�$^a�/��/�`C=���#�H�p׻dr�D�O�Q���r��l	kb ���l<���qw�3�o_�|q#��3�p�nn�cQ�[����;#�ZO	-u���|z���FC2\�4��юK���Li&JS���І����<�E�Nӊ�Y�SZ�C�c���a�P3�n��C<��zv^����t��r�Veck��+�֬���������WJa����fJ���.A���g�S�p�t�}@uZN�;���@��l��	��s���#���[�O�Hx���9������P�L�a%C��ƽ~E7�-[��Z�K^c�����9�h�2���^�t<�{���q��-y���w�bbb��7�[�4m.�N �_�l_�O���2�z$����о�(��,�9ɮ;`&�a��i4|�Z(�W��4#�|�f55���0�L_,���l�~�)�	rE���áM>���:JX��*�K���O�$�m��݅-���zc�t�up�á^����bw�9��:��Ա��"���Ǿ�/dEG~{|�6�t�K���}��M^o�5ؑ7{؋�}��������v��<�u&˩�CF;���>�t���(@�3���%+n�N�xN�9�-�/��4��h>�6a(Ub���#��3����9��b�/A[M��x�� E���m�v����xХ�"��U��������^�\���>�X�(���X9�I�����y
�$BL��iџ � �c��j���H�4�-^���,}�(�ALI�}p��J=�ܴ��X!��Ւ��vׇsj%�X=FJ�&����2��d�-.�2pӯ3U+�~"f�M���s��e�nF9�����~~ѽ�ˌ��V֛H�*�2�5Ϣ�����z��F�K�v�O�Rd����l��2'/�uN�6�"�u܇�e��å|�h|���aCIT�{Ph�ie��4������-	����ν�ΊE�I+�#���g�sL���ZW}��n��iA=P�!�R�Je�/�����tb�-é��8lo���r�j�Ղ��M���6"`�äF�F�^�fV�h?�.��ɺ]��-����$�0�6��|�ڭ�;w�^}�[��Ɩ�)��T�V�������#�^���S��jÏ�%Z9�n�y�G�G�����=h�:����Ci���G��hQ�
��4W3b���䥲���Ӣ�"g.��3^߹���H��ݸo2	��-�a����qZ4��X�-���ؿ���ɨ��S��(��4��ϕ���T�G�8W~U�>�Q5���:.���
��|S|�4����ԫdȩs������;�GؿnZ�]��6[����šS-�Y�޽���d߻��DIW=���h��2��2� )����)ޠ��E�Ļ���RVuH�/��v9�Zވ��Ϣ�y#�o�B � #{��ѽ4��@�4h7X5K։O�2�US�_{�N֗��h��� �ʀH����q����*�(ӬLM�<��ʹ]t�E��Z�/@@j�\�a�	���u�0���g���(��>���xJ;z�����K�-A�D�n�,�;Cb�Y���@���'�����w_�.�YL?��$�[	 ^y�����g���9�<�*J�&��]�xvh�_���n���1�-�AԤ�m㟋ܪ���+#�뜊»��� O{n�6e�V3��n�Y���Q�&�$__<��$��ɈT��s��;Kݶ����1^�phJ�\�*^O�50�=��l�+����3�9�JW�"�2�����Y�R�@6�<��f�5��`�P�[�Q�)3�Z��,�?4�C^�S�Uԇ/��;�#/��^3�&/���[�L��qlާ$�kJ$!���}q^
m����s̳g�#��u��P�0h� |CIԚ@��!t4	���MaN�=�	˗�"%�Q���d��\���ѫ�Ɓs�/q��\:F������������ L��)�g��?+�^�=-�(�n����������\��p����]�<R� ���=����|^	~C��(����ϓ���4v��4Y���~��`���:w2mm��������f~ˠ�Nc+�rK�������A{a $� �n�7�P��^(��3*[��X�_�P,�𪲋Lq��'��(W;��8���###�j��뀛u̗�qŷ����e|�@�����:ؓG.�-���p��{�Dv������J;ߧ���O��z�ì�JC���H��χ�n�{���������
�m��C*6��Q�ٿ�i�C�
`��v�F�s֖`��&'�+k�U$fp�n�N�˯i�[���uW��"��u��	 �\�$Ch������^��(Q2���
 VW�� 5C�ػ[�?�Wf�W���㌕�=����].�P����Bw����>Hk}9�8�˛.��(�ڢ*�����S�l0U����7��,����N�t ͂鈸ǝ��sӟt�ܵ!,.*�����c��y�l㕟�n�m%m�od:�$B��I��{/��P�8�e�tdv�e�?����)8��ioj��@��8����+�2��﵋7��ħ�>�i.�
_,���+�07H240��Li&�ĝ���9n}Z]��*�>-�:��E���?�'�T�t�^����lM�3\ur6�A�=4��i4�_Un���u�@�)	�|����2�u[_;D�3�$���jhh|��;T�bׁ1�sW�N�s��p�ys-��8�y0�ǫw�~(/�B���S���a�ȣ�����o]�i�FHꓴ��W��7�`�}_��fLi�Z@�d��d<�sw?IF��dkD	�$�$�,\�o1�_RRb�D*���[	�}�����r�wi)��}�d�������Ŕi��#�]6���A���D&�d����&��Du���*���}m��^"][����G�jUt��[U�3�E����>��+�D��u]}"\�q���'��T][��N�������V^'\�Ƚn�cw �G`�8�d�Ɨ_��7�ׁ���2��%6��3'��j��W8AAP>�M�V�M� JG�	ԐV�=9����CnFYS�r�H�Rs�h�c�ߝq�R��>�h��hf��'̓=���}ig3�M��Q�["{7��y���`䆉�V��q�z�h�iAAMvas8��L\T�Mζ7�T��Jr���wC�(1���yO��;r�8ԫ������g�}�کҁ�"&��EZ�
��W���a���x �����rTO�R=���i�Y�$**�I�<�1E�)፦��l��/t�8��������<�L�/E]��c\�>_�.����<�����@<Q�\�-(++PGwA%�r�}+�a�{�2"�~|�᧔��|���)L
�݊LȚt�� �o�)V���^�����'��+	㹟/���>7ޔ{X7ox
sga[��~�	���i��D;��H�H*N�Z���N9��$�$� ���n\lb֏�}�k��I-�`V������"#M�*�BG��;��Oˮd/�2f$S�4����VyCw`Ǎ$b��$��=�>�/(�v6�{Z���D)[-
��LX�' U{:����|��`���k�S����8�31����S�U����,ҿ���:�9�����jF�W/|�T���M�4a���+(~ɪe%Z��ObF"��b��1�}]I�f�ܤZr�%a���TK	9�Q-i2yZ��rDE;��������)����ȰQ�p#.�݉�V(S������3ׂ�gftƱfy?N�G2^�%�$WQM��U�+����ڣ����2�ll�p��|Kt��s�����!� (��yaW�|wx|�M��8�Ş�'��΁���# *9��&�u�<�n�s��eS�����ִ��_�����i�z���ܯ#c����[�>�wx����BW�.S�>�_S#��(��Mr�p�7ӺmL��������3y�/��P�,��0e����T��b0���F��x���FEə���%IQ?��kj_�t���[��q)
��Ǜ���0�!����2}�x���������.#���}7����L)�t �橲�D���z�e�*��~�t�z���m�q�RV�`��R x���	��n���޵r)5xQU�4���tFM�=6������� �*������e�#s���etO0qW¯����0W�N���s�F�4M�8�no��<���(��KG��i�����_G�<�Eݨ)��e-A�v�ժ���[��e��iߙ`��$����\�L�;���|�	(� z�,�e�t�ܼüE"����1qW�vk��rM�7'��9�>8�����j��ER�\ܴ�L6#�=㌌�M�C7s��e�N�'�68��2S��:v��1�PY����~�qR���z�Ś���w�:lo��Om�&-138O�͗Q�|�+.X���!n��'N���Æ�m�.��r�"�w���5J����Q���*1ʴ�FiMB�ܒd���������R���T��L/7��\�f�x6���,�����0?�fV��7ki'��64RB$R���j~��3��}L'�	��z6�0������Ŋ��=���Z�1��V�Lo���Vo�	��T�QI��3�:�����ǜu'=~݆9IތK@�����g��O������G�fF�%���mn'����.q��u;$|���%Y$R�z�U1p?ш��2 t|��k�l�c�%UP���~-p�@z�Y���ޓK��d$�ä�[�]E�F���I�4��|KN��b^�5�pr��8lܜ�S������d�[�6���h��,P|x�9��" a����.L�V�rA�[d���1��-d���#<"%��B%�;�YB�79�7�틗|��-!x����t�
����Z��f�Ĺ�J�t��@��~\9�K_=��D�!6����,���^��ɿ�CU���������a�������LZ�d?_�6B������Vyt���-�}5����%���?�ޞ���w�
�j#��NU�������9{��ը&M�\$>��XU��q�z������VfliO��Y�}�
�"%�yh\�94�m�ܝU�u^��.x����$��l{����C����:4g~:X��AS�
p�D�����!��!/�~qeL�Q�K`���=�l�vEZ�<��J�<?X֓G@��/s9�z�u�d�C��F����O��b͹ �Qyy�ϋ��&w���/�`�ײ�����2*^�(�BϤM�����!pU��=h�\��p�$5wc�n���5��B�e�+|�g��^�k&q���jn��l�x0����.���ۘ� ���Gr�|Ps$�a�P�S/���H�������j��o8w�����k�
<������������Ё�'6ǵ#ۭb5�-��<�A���{����N��Ӻ�������TkK(��u��3T�~�[_,1�5����S�$��k����&ey�(`9���k̠A�6�W���Y*�g�9l��Lv�8�}�3�+�Di!<�#�k��	[�u�c��VWB7���5������o�`A�]
�c����n��rCo�![��֏�����GF)�A�{Mڥ�l4���c����L}gL篴B�	ߒ�s7}�z.��ඏ�%[�h�xu5�u@jI��ZB����3�[TF�{�S�Fܦ�R>5i��,��B÷A��I�0糨�襬��4�^Vf�R	`�#}�����hþ������������W��Y�����ͦ%5�邷y�G	�N�_REέ��X:���а�4>�[�V��H�T����^M�B�����tG�+���=�o�:�kx��d�G���,xf�={��+P��{q[�<��m��/�u2�����6:/�F	!F;�؂Z��}�1�z���#Lo1]:{�А��[�F ��]ē�
|+6�S���L�yH���h
�Y䮜f�z�O�.:Q���0��^䪓��p�)s)
��z ���OZ'r`)~zz,-G�R�ü��C��jQ5�tx�f����.N�f�����,�n�ޒ�p�!0���ۏ?�neHY����.A8�0�+H3H]��^�wٝ�p�:�o�,i�^!]�_��*������v��S��0�)���~���Z����bO�uY�����_��
YCi����0�
G��Q`�� `/|Գ�T��i#�pUKvR�u�ִ�s#��2���S!����2_���1ZϬ�'���t�͚<�{���!���@W�$���@H�+;C�ZRq���I�4]��s��3��o��.�#����b�S_W����9�Xjɞ�Ў��=5�I�*��[��^���8�t"8l)N���Wo����!BH��<y\����q�s�T �Ц���cV���?���7��Wri����~�A�s�
�g����b����ka0e߾UJvov��^w�����A4�a4�t[�0��9h'��"��R�,��?�MP&Y�X�41�G"��D��p��gr�S����F�ԭ���O��WM�`c��8�J�yɤ�qC?��F�d2���%U)��S՝W��T{1�Q�,���R���瑖�\��w�B���H�,��]��O2Z���ӌ8=��&)���%�^ ���j�✃>g4t�9Q6Y�����R�PU�ڑ#�JkSj���z$9I6M��û"�&HuԜL"N5�(d�hN2X	�v�R(R:)]|�h�c��[�/|������W���RUmg���y��ꮜ�H��R��Vj�YN&�:��2ԣe�����+xO�Z���� 1v_�N<Ɵ�M��-�t���a�IPr�ƾUڄ�;�(���ay�9��S�A����i8���.�I�x�>��O���$H������a��y�JLIq����t+-�p�Ǿ�~��2
����ڣ��Io�v#7�*�ڗ���W�����;�Jj�����0_�YI��~$�e0������/�Q�A��1���lF�c_���[��V�3�<,�z(���V��.��� ����cKB���Y����C���i�R�+FU��]|�z�=>Qb������++5��2<�3f�+�g�T��x�+�@��d��f ��y���6�u�lS���������
`�4ȫz˿.H��7�#��[yG�����)���h]O�H�'��s5��ݯ�R����mΤ���ߒ�j2��&/�#�`����Z=�M?2��r��&$���ۓ�ƫ5&5�a���9F�ժ1e�����C�굲�|@R(fЫ0��,c� �9(w�L�R'�3��~��3���I�$g�����</�^��`��k�Lv6���U�mv��#�tȾ�a�-\����/}Ey����/���_�Z�f؋n�7��/1	�^�^>RrL,�M!��&AN�3�6r���n��< 5�@�<�#hB^����=QO}�58}�����]��MCJKl->�ѪA^:�L����v����C`�7WPkK� #fqfi����?�c�����U�����[]�+(�h�!�����hﱦ��{�%s�Bb��)�O�(�������}�rrDHU��Q�=� ��P��w��(�H����'�z
������QK�^��=�&�ˤS��oI�C������O���!�w�����S�p�eF<�,d�1��CmاF�]n1���8꒿�0e����&����y	��n_��̃�B��I��c���
���S`�}��th�Y�E�X�ߣT��
]���p��b�P41B'2�0I���q���H�Q��Ã8��q3��N)�/��?�ƴՉ&C"�0�}�}�RH�#\�cA�BLv�ӳ!��Q'�T���bd<�G0q��o�Q�H'w�2j��D���gq�#��f
!վ�������< !B'��X�^.���]��@i�s�R�T�T�`���?@a$p�&�{��%���r��F<y��w�GcI��?" �����{ �D{�|7P�%��bo�|�0T�������
\���qE����}���ەw�UN�!�����O
$�yF�MX������cX������ILtb��5l�xjDzB��n�˟�@Mf��hZ�dy��t��١�8P`��-�J��Eޙ��e�S�w¢����A"�o�Php���v+��f��9�D�Վ}vmuP��Vz�Y��L�oR��+��0�e��;S��)������-s8cd�j̀��+��J�̷ޙ1^���	�\��L�}R2a��
��&ױ1l먺��_��D��8B�pE�sy[k�)Ӥ�Γm�Fԟe�ۍ��9��֑�(|^M�K�L��T���C	\���P������E]d�Z"���SzW�����2�ʎ� n� �W�|��^H��A�[kq`��|�+��$��ÿJ�cEH/��&o������(CK3�P�����5
)���Cܤ�G��[R**��M�BJ�r��$)4�
�!n�S#/A9���|�]=�*�R3�p���	V��iׯ��,��n3�� �)�(:%���w"��)5��?�{�^�ʮ��q��7S�V�j-���yYVN�Le�#�ǴY�!,�  ���IDT��}C�ܫ}K6�bh�X���N]čE��\��܆�=���Sc��Z��[n('q*�P����.��S#è=�#�\}$vm�
;~�߰���,x{griE�3=���x(�Ì�E�&����F�������#��׿���f�2���~�a.�RZn�Iڧ�zHP���'��bDו��8��X����X�0�^�Z���J�}�y��"Ⓠ@R��
�/;��>��hG�rGt
l�Z3IC�|Kl`���� e�RXg�)D �8 ��`�sO9�q�h�)�X�i���l1�5X�(�@��w�5,=5|y|�`AUF�4�r}�}P�iFxN��2W��ϱ蜘\�M����7G��pȞ���J�'�Ӄ�;%C7�"S΢�Q�J���r�n�� 3�-'�O�}����Oi��/j���������|s��lP6���yϥo�-������O���Z�d�-7���rǥ֍~��SNRK�Zo6\�$���ͼ=�(ǽ����m�.B���r�����̮��d�S?�����+k��|�����/ܫ���������	�o	Ac��%������ߒ�[��oKV��\�u�����[�K�߼$܇���h�E/��f�����IrG8Z5\���0�cN���\t���tUc x_�^�޿ ��$�˿�ﱳH�K�Z#'4����f���c~�~���RV����i���Yh���+�R���1����k�W���u���"�����gH?m�W�C���Ǚ1�s�(������߭��-��%����KR-���ѩ\�u5¢k`���@�>���'R!,�Q@����YP���њ1��;�ەR��}j<"��e
��>9AF���|�܅��$3Bz[�B"��)�틛q��A�Z-�"�q#yv>Ya��0"_OB#��](�G$�+��y��݇�D���{�~/�
�D=�4@f�9QJ$��@YdO����2�<�u�;����k��rk7��P"e�/�GK<cq�
��i���,���ػmV��k�,㫒��� �{�t�g�L��4���d+8�
�J����U�	�&��d�޶��5Kʝ˅� ��E��(Y�CuX��Y�_�(�o$��2��"B"J�������c�����a��nKC$�c��s�r�I�Kτ��.r����=w����rf���W�{yv�x�^<l~X�j4?����'B��}��+�(e�9yzh~3�~rA1���k��t��k�����P�C�/+��w#:gZP�6o�g�1�b�g��~�sG���f�y���F:;��E�
��6���]��bQ8�ި3�1�Qzܾ{�KN��y��1����Ì���V���գ�t��\QK1�����}�ۛШ|�T���}��q>��r���0������AK{����Ծճ�5x�MVv��:�U�a�MӼ�H��>��T�NOө��K7�k��5+{}��p���q���Ƀ��%�:�j�����o!�����E�j��K��0����|�Ϣ��3����Va�qW�m�wЩ!�q��.=Fu݈ʿFk͌\����=���9ꨆ�y�V��%=��7�����u=uؗ�LW��X+UO8�'�2�좄���߅`��֬���r�	^�Ȏ2���>xƟ�������gFN�^��h[*�X9�	ƶ:d���b��[�h����rR�ћ�6�\=�P4΋��	f4rr�dn��.03r������;�&5�ET�7�!����䌰�*�st�_���
,����� �����^)��k����z��iSu������ �.���/,sLn~Q��o��^1�ߤ(�����Xspf���1ܩ;�hC�<�c���dq��r¥0��0���9;�c���`�%���e� �+�_��|��u8������}2�8N���צ��H�]��F[����BX.	���.>#�zQay���c��t츞w`쓻r���d��5SNο��UZ��O�h�Qy
��|S�Rl��9���3�������^O��6��$
-�����lGTa�}��i����].s�߉�Z�AJ��9꼍���:.U�� ���+pݻ��rM�{�*�QO�����/�*pU���4��wtP�ӳ�0���~�[Y���|�G�K�G�NO�fr�O|}�u�R�/�N�+��
�󽥁��{L�U>9�n:]��פ:6��V �����BӮ��촏����g��� Z�`bF0�yT�F�DӍ����k��5`�P��ܕ�_�\S�h%����R��O*������1\�AT�'��\����5ٙ� �$��_�r�|ȑ
��s���G�3��<�U#9�NW�W0X}����L�O��E(p]��/}�a���F���CQ�,l7�����T��3W��%h\p�É���H oA% ���6�}`��k�@�5.D�F�%�\m8/���{O���ꝧm��)k9 �0Ό3#�!�<8aZ�����h�,|,|Wn��8��F�2*�O2�-Sop��Y��9�-����M�����t!��0(���ԛ�r\����������������}{�O#AD|�׀G���`.��m�əC�XMH�5=�:���.{1���VT�q�e�}x���.���3��n��Y�P�Uф�w�!4o��kF��zQ�,u3_i�z]w|���1]��M�0�5�퍫�I\v��T�u��(��v2�Mk|�k��������g+��!�F�z_Ttz�b7L�S�8$�����a�7���/*������X��7}1���d��K�[<%n�-t^�yrC)FV�c�#�����a.D쏳���H#�����h��؛X
�s��,J�v��Ub�u	hc�~��*���K��a������{�}n�)D.�zڿD��=c��$i?�Lm�Ҡ��i�9���y���_�ĵ
C��Qa8�wt��]F��٫��qJ.����]���91����&r�]%�u����oYt���E�b���*��k��r+��y�z^+ϻX�w,�c�.��9���^ɲ��[gր68��gW���1;�`�Sv�v�%�:U����A��ŕ���ޏ1>֮0�,��E�[BM���(�����e��� G�{;�w�"�}C���H���4�CR�*���=�i�z�u��mr����yH��R�(�@bI�p=�����	t�B��������zr �I��c:��gɯ���%��K��\4j�yi�������J����x;���J���1�������tvJ)q{�"�P5�J���f���nخ�%����t�pr׿��lN�7 I�ïI��_p�9}o�+Y�r#��;$ꞔ�G�?!$�xRC���{F]k�d�u�{�T��]/�t�"�ުyC�*����.��v��?���P�q{��U�J��)�h}c�<�����Z�����N04�y�ȹ���p��7��"��Ɂ�
�g^�m�̈́eO�)؍u:���UM�s��K�춠 ��uU.���qIӻ�8{9���U��ׅ	>����?=���i"�o_����-��l�6�(.=���|�j�_Pk�\��
��1���h����}<�6�+B��_;ЉM�b�Ud+]����À?�LU�����\r۠Yxa���/m����n�ױ�U�Vs������JyL�`�l�jZ��YGk�#�3C�Ʒ�%��2�{-���R,��F"�U�Pݽ)a�8�"�;].��{rh�b�O_^�q�V���^� ��G̪�Rī�^*k�0跌k��V�*H&{��A>�T���Q1�v8]�'s�
 �au	������%��t�<zߜH{�H������qK�����$5{�ٹ�U���e����ob^F�:p$Y�D�q���ԗ�OH_\�a*\cz�.� N�R|Vp�_��j�w��N߈3>��.��11�%y�*�3�(ް�n�au�����+gޝ��bY�t9t�"�M̑L7'2�C�]���t3����H����feL� 	 [~��N�='�>=������J�c	򀝲�o�bD,����rsS$o�@Ec�Th���-}x��X�,շ�,`��U� 7��W���Vc珩Az_��������<*|���!Jhd��q2�>�������7L���y�j�;~�4୑DCw`�af`f-��[�	���f�0%3�	o$��}R�gs��)s�d�K�V�w��UԮVbP��t^i�L�b!�,P�j���ŕi��u֊��QFY	�	j36b��t�<uddߠz���:)��:����J�@SkE����P��R"T`��V=P������-qfw�����-'������ǧ�߲�A+�#m�g�1W�3�{I��a�����G@6s/H��О�TM�T�y,0^�X�Y�5C��ɮ]�д�4y/Q��, ��1����k�/�4��+�j@�٥�o>pW(U��I�{3/����w������Z�^S��.�x®Dy�W�{_��
F��B��=*i}˪�@m��������]�Ղ`���u��ӛ��V���*��GG���gIʹ�+��j��T��G�P&�Yd�`�n�;�zX}��Pt�,�kH���V�M�}��ƃ��6��o�2�l.�< �IP��<���QP��W�����)J�;��v kέ��J�矮�n�&�d�'*i�B���Y�5킁�ݺ�#I�cM1D3SX�W���P�ǀ�����9�XB>�����R&� �����MC�+� �	�B�U���p����mU?��|����;�������?}����g̱ĩ
�ڌ�LvدΔ��f8͓��GB6����.�4'�0�"����pNq~0R���9�s)�|��W����j�^~�y���J�;>},�o�u�2��%��$?�z��d5_��f�
�Ͽ1Q�A�7p���� E���R�RϷ;�'%Y�{D��6Z|�;�� *�Y�E�7p˵&=�yj��QqT� ~�;��+���?F{N�sb���y���s�e��s�A�ʑ��"$�2��G@�P\�&�[yd���H�.��� gٻjj�Ã�V�}au�*1�B����3х� ������c�3<v���������ڰ���[7n�]8��!:����=Vd�L!3]�Yc�����;i�j��͡L~��%����(-Su?��ݧlL6�'�9�G�9h��>�����n66��|���������N'�78]���xf�F��s�R��n�2�ۈ��эd��՚�=р�xmo��:�K0� "?/�l>S�j|g�Kz�T¿�ac��oczP`�[�'�m|+Y�m-��"� ��bTd�H`�_22ͱ�~!�6�����7N ���	�`������T=�,==���M~R�0uێ��M��$zٰ������bb���mXz�\�o���f��El>��J�\�?S�=x�oK~��Z���x�#����6�V�ؚ��51.�����ιC��A��������.�)pi��U�'$^��Z�qǃ��4�l�*��e��$ef挭5*fA���K빽Y�!��R5��eF1�
�#Û� �(G=}��]���EO0&���k'W���f>������üD�� ��+"<�Y�r�� }�=ui!�p�K�S�M �0T���VH��#��C�����.̣�#�.e��
�Ĥ0��x�[7-N:�]؃Z1W`޾���݊��pۜ�S'?��:ٝM6�0}dR��b��6�_wP��Rz�P��>K�7L0'�A�����
����eeC����H�랁�马[��C�����P�͉43�w�� �W�ܻ��8��I�uW�%�i��"���i��
��ײ�h�����,x�Op7�d�%N:���j�jK%p�;�ax#�1���z+gsDd4�7Y�}Q>��n�vO�����j=
"'����XC/��n]� �@�+/���<�8�Q�4�)�g_��Y3��6����@��u��OE�1�l����ǥw������Tŭ�l��5�ە}�OHE$��%�O� {�?y&���zΫH�����:�R��E����ˏ<Q�(�9�3��I�:��ˊ\v*��{|)W�5�����t4�7I)�Q@ȇ�j�;���\�~�|�R+�����d��.����k4���}\�:v�+8Xq�1��B���˯�����n��"�wn�q�"1װ�H�3�Upӛ>�����FT�8�Bj*W=�55���irM��,�iY�o�V�p>��!b�����o�fB��3��`{^��*�Q?p�
���GZ|�Y������O�&�<q�u7g��$P(�!,���Bٯ�E?#{����-�	D� �Kj ���	uu/�nĻ�	+r��5$S�@��o���p;��y�٤��4?���HX[� �iwķ�q���R�]���@�X��w��<�#IrE�k-3����	�kLҠ� lx������S�zX[�/UG/G����:�P	Е�f"��s��~C�-�6o��B��1ٱe�l�vVSK�'�-2ڒX�R���:�7���\r��T�#��Y��뷞̑���ke���V�WD/��ڑ��,tw���/@�4m�\oJ���A���ܳ"~�����'��I�TGc#�b˽l�0�〦f@�˷�Wm���c�X5�-��x6����Aէj5w�ݙ���7���=Z,(S�k���pī�ϗ�?��S\(Sz�?�*PD�ޡ�H���V�&�?'��A�砄T�B�X��X����Uw.3�eYU,���XnV�r+�*��bR��U��z��Q��C�f� 4��X������}C����ؤgFn��߯+�H=��yf���DN�2�������:�,�~5��A6&���I��-�1��iա�I6�^Vϟ�Ome�����y�h!Z�@�-�ݾ�E��:ۓ�W�bu'#A_�y���U�pgn8�~L�Syv&ij�
C��{eB��a�[�vї�>$G>(%����*镘�@QR�*�����|c�)��� 	�[Z���(�g<%�v1�Ck��H������b��/�ͬՃġ�6�Pf5X�9�"���FK(G��#�+ŕg���O�ԍ���rǯ���f��R��嶞L�r�D
'�&dbv�c|�fE��j�f�Ǐ��^�J1Yx�oU�2yq�U��v��%���>��g���z|��0E,Nus�@�l��i� ףJ�͡��n�߬��/�|�?9ɬ�f�\�� ���U'�X٥�zY���}��MzK��ww���F�@��pI��Xt��rr�~��Ũ`�'w,�bU�v��x� +K�TL/�"�g5O�8��i�E��|�c<ŧQ�����7<�Kc#�/ �.D����6����%YEY������V���7���wCG��H-�kx��,V���$4����2Q�Brh;�
���{�`�@ ���Vbf�<��ʿ�d��Zs?��b�l#�4�#O������B�'���v����u٘��Ju=�6����*�w/�Yn/�����}r��zϻ�?��P�'i�ýc�~�������e�q{%u32�|����{Y^���Yf|���Ѭ!���b��l+XWǡ�f��m1O��k��J��I~����ĳ}
X��A[��o-��_Y� ��U�YC�^��jSA�n���6�_#�`"[Q�Zz�Q���f`�^݈~���Y�8@��@8���� q�M��k��Ўw�C:k���oI%�><��Κ����|ںYZ�w�/CH�8��=�fW�� �2-������}�ֽ��;�+}#B���w/ �d��� U��L1��u��T��U�B�'-���֭0��Q��H�m�g%��)��o��l���t��H�� ����W�L��[��j�\h��Ԟn)���7)Ș�v�l���8|]�4�o�"o������H�cn���0I�'{<�TN�:��+n�d� �*��qxU���;PًsOo���ж<L� �B��s���s�O�'����X�-5���*]�;8���)�'$�E?�y�U%<���*w�l��0�������T����7b%yP3��2IZfu'��*��@���X�-���36�Xa�i�<�r�4N�2��e���Zë�c��E�ɠ�[�[1�q�*�\9L(�>��afnJ�3K��~��[gߝ�jJ� ^�����#�>1��~��vYH�����hc�سF�� �ֈ����@t>k���lz�\r�҈�ҵ�z�=l�~��JZ�r����D̈Zxm<d���H�Z�Wg�*��g̞��O���ybw��������S� U�M?��0�af%�FOݛ/B~�2,/L���z��u�!��s̭�{��e�)~+�M��i
��dC�qqr��Ad��wD�J������m5�O�9ɹr%N+Z&�Y+z铜�s:�0�}%��ɶ5 I����H*i/	`,.�,7��T�g�@,�A���T�<�흹d�y�RA鎂����� 4��7SAC��!�.Tօ���
^��Ⱦ��WI���{G�zBM`EɆh\x�����@&u75V]���>�ȩ��p-|���x�49[PN����/��Ts�t��}*o\�LJ�Uȿ�T��Z�61#�.�)'w��i����s�ŷ�fg
8]C�T�����E�^ m����i�#�׽:ץ>ίTb������ｭ�L_8��r�X���(���s-k��l}26��f�/�W:�"��e�xɤ�DUL��x�����[FEٵaÄ�����AI*](���"��t#݈*��("�=���0�Н�Cw3�����������Z�Z2׎3��8��s���IQ2> Z=V2؃���X?�����t;�)KF�:�w�>E:BU�vL��_R�'d��ӚJ-�1R.���M��L�ӷ&Oqmk�N�Ɋ���Fc���dOέ爖̡h�(«?�P�A��IQ���Z����d�ݍ����[�#KYi6jj!�|`�f�R�F�ez+�}�E��� DW��ƭj��vp)�*�tOU?��j�=W��_��}��Lu�l�]�X��O]g��t-^lfO�N�o�x�d��MU��%���g5@��P���}+ޒ�x-�&�0>���8�K�{/��	#n�m�ۛb��:>f;�����4�Z���_<ʞм�x7��2s")�������D�z�FN�iqN�AVz��3����-�IQأX��� �=jEIn@��|�n����|�]鎀�����&Hg�-�,�>ձ@��I_��O��/�w$�!��m�R����q�����d�b�n�D�g<r's���y������,_�}ձ�M�
C =@Y��ȕ�6�z�c�o8/���?$����'3!���Ɵ��1oH |Q-�>�����<�6�6�j�5��J�k���r��o�)���\- Xy����p�&�P͕Qeh�L�y���4���.�� Z���Dg��mʌ��!��YЪ�����L�� ��Ð<�zh��P��#��@3����O��:K1���q�ly�fu�>бF�� ��1���_"��jgi#������O���o�\��r��V�ǜ��+@+�D8ʫ���x9�^>k�Q���8D�w���H�r^�{E��B?3��Ǵ���L����!�h�S�����Q�,���胖)��Ǯ�]+�6|Y^���71�Y>���[�1�u|-i:�vDf� ��q"*���c�P�\Ql���z���;!Q�g�36���M���i9�m�ꁘ,��ae��;ic �M�����<a�n�5PXCK��^"_�Mۚi
p!�,j����?~�vJ��S6�4�����ft���6?#J2�P ��ș��}׈�Pi����iZH6������4�����3��B�A�_��X&��Tq����d<gw���*m�M��N���D���ͺD
���==�$C_�_�]��Ǯ��;#�d��d�B(�']*t��:�v�O.�I�I���l+h��V�Lv������e��Q�b�ݦ|�,c�q���5�X���phY���Pf�&�莻�8B��r�]��^� �m�.�B�5�p��ĥ+��GI�MaHn|�t��x�`Ո��ㅛ"�,ݕ��̠�s�nׁ.��	%KdeE�yc߯򲅠�Zm�2��Ko�c����������`O��C*� ��{jߒ�x��$�8	G�E�ɜ�>�w�av%AΞ݄��'ޑ����+@@a�� ;�U����:%�%/�S�	_����[�-�y[ջ�ژA������k:t�:��č`(����s�!�-)���%�f��c�(��@��c�Q��WЊ�j���N����e,�ui��օ_�n��;fM���)�طdWbPlS�����Xd�H4!��ES��g���W@(^��ͽ#�'E�Xܷ"w�����	h�wbي�6��y|�6�s�<���F�u��1�+���H!)�������J��|�����9���ꮯ�钭w���/y��K�O��	�Y�B� }8������o������(�/��?
[��vc��r�m�}�Erһ��z���l*���`, Ѳ�E2ڔƲG�~cs��V���>!e�� �'��<^n�kCS[��^��iY�]��#�W�"����*��5l��0!/��F�cS�R������U�����m�wA^E������j��;7hŴ���)�A׹�{�~�Gȩ,ym����Q�n�>p�����Pq�3��r5�MR,�{��׮`�$iDY]�m>��ļ����%	����W��Dlr|�V�$����CE��y���p�<Y����ţ�E��;��w{�	��E�[
E�s��D���uΎv3S ��[c�#=�IQ�q��C����!N݇Ib��X�ݟ�7�=�9�o�*�m�S���iΦDU��?H{����2Bk�ˍ�%� ���):`�r���Ꮘ��oԇ^7^�+i�C񀇨?0#�\�j,�8��IVs�A- i_��R�Φ�fx�xu,�Ci���ڛ�8m=u��hޛ_��r��C�X�s��c���#޳��fzRѽɶ4B�-�~�y�XO ��5oU\��*Qf�N��z�ދ����H�ԕ;�Dծ.�n��&k�@��4�O�l/��7`�/�s�6���im4��� %�|ӿ[n.��U/����]�_�f��e\=����ͲR���5��@����Q6kh��\০�������謿,ګ��P��s��������V7�Ϸ&g�~�����Zx�")j?f]�˝�P��-�n��ii(h]��<��$���kł�����ٟqJ������nc�j֞sr��ç�Vf3���_�Viz&�����~/���-�������"��
��n���7u����ߝ^�9�������!SU�k�����밷���y��+\���*��ƙ�^9�x*뜆�y������Q�ܰ�٢�ڃ�ƥ�ڳgOA�$zxt��`�j����#�<���)���*��������{}_!�5����,�����!]��F�b��Β�B�f?Z�{�i�H�i�ڜS��<NN������Z	�7���]P�NW)������K��}�{G6��Wd���D)Boy(F�o����v�}����g1�m�r�'����s�*��������)c�5<PcWg(���W��Q�����a5��N28���p�L�I����0����I�Ĵ��TӾEvў��~	�������n�c���#�X�Ï��SL��5�k�����K��J@F�y�����FBH�}����G��␻�cO���zv�SkQ'KK�Ҳ��5�iÙ>��a���d�y��B�r!�O���]��"���є���l�X���~7�eP)�s�J����fz�']^�S
ЮCُ���sY���
�`jSɬ���*-o�5���؏�5y�3�"�̬FjJw�;Rj;s�WJ_�Nˬ�V��M� �͗C��	�
�ƟB~�k���7I�|��(�A�� ��C 9"<����x�sA�ׄ4���~4��iيRn蘏�	�����j�}[L� ��¨ާ݅~�dBZ�9�f<��ߺ�U[�裱���6��С�IR��g<Eǟ�I�<wB�ȼ��Z��lO�]mR
���q�a�%�'�w��ufS�(A���fݪk%�t�(Rw��o�h�3��,�U]��ᘢ��b~O�/�V�9x9�!��7��n�f�ބ*{"�md�Ǿg�&�j����'L	_�:Xsߕ֏��9��)�'���j̍�aւ��J����N�?{y���5}0#�X~�Һ\�����Ҩ����j=H����	�)�Cg�@�}b�J�S�~�*QZ+�]��Ѝ��gIѠ���w�����JV�ܳ�>>6����m�Z�@����<�d�' ��ZL�0b%:vl'M���ߛ%3�5U }x<��V��qh�
��ݬ�VMh���(�2Izq���ʪ����b2��B��p��hkF���r��2���%�	7tPa�j�:sb؝7�Y�8H��K�c���i\���GǙ��V�\n�u�����a�9(�O1��҉���]����m����!4�ڭpn� ���O^�z�*Z�7;6�{��Eg�|���.�6z�	��8͕����d0�՟5�\/�� _M��,�? ��Yta�:�����6���ʠV��:Ir��
fc�*""Ƅ����t����ϐ����EN�z�{���ǐz�mߤǭ��Ж��� sk�^���Iq��0sb�v@�m�o�$�CDC��)A�c��3]�A�)zA47@B���yي$��>['e�ޚv��j̞"��s�_M�T�NH�w�o�ۓ83jt��n×��F�<�JN(�,�p�,��"!^Kz�[�Z1�y��`yz��N�_M>�1�4��'��s�,VتtA{[�b�(�-�a�{n�V:�C��{�ʼfh"����u@<���h~�(x֣|����������y�"' _Dk"�2<��q78_(�xb|b �e?hŢ�X#!aQ��O�艪��.���F�I�/4W�$�n�}��4��>�0��1PFJt�O���?����b,��y\_d^�����Ƒ<<�Z�-5˜8(L�,���w�b�'��_������I��"�N]2ҡ߰��>|��O! >K�t4iyfs葽�b�f�IzF;#i�:��U^�t��XUpݪ�K[�G�L�C�|A�%���Q��u��5�3�Q������˨tNF���\i�����^�����|��}��Y'a�Xb/	|m[V��<���W 
��"�K����ڍ1�V1�P^L�����8�N��;�.�h���W5�i�kQ�J�x	�Ј�����.�SUa��Ec_���D�T���!����9�Oj`��)�!e��z�`����8��,�������TA!̜�B#m�}��{�������k�zƁS'�mH��n�^R�g=�U�M2�9x�+��,H��V0pm�4�l˧���մI+��l41���#�Ϛf�-���O�k�7��5����:V���1�3�	�C�Ɲ��� �A��Q �U�W�n^ή[�ێ�8�ɿ�VP���$���yhh��CL,ګRޱ��.�9qYR��U�ؔ�X��9��-8���|e���O�f��D{�B[�5�gEG"O�U�F�H�gg��*=-y��<�嵯��Ë�@�֭ ��תH`�],�*��CB���s�L;k��cv�"Z��;�+�I���C�����╾��^��|��o���W3]���k2�+����7189�܏�U�ojF�M��ߴ�X\�$$~H�`�J��cR7�)v�2.ǯ���͕�������{�>ᠸL�ȫ��TI���e���X������m}-?#B/!��(��"�t�"M9�S�N˩����ֹ'�8�I_S.*�FB����h�K���nV��_KR�����z���!��%�Y�����t����?�tM���]2H�9S�}.M���t1 �s���\�\=m��R=�g�����=��O�����]:�A�[��Y[W��������'y kB���Q���������=�Y��#%�]g*�i���߇�N��M/Ul��?�c����H?�8�s���s����G�/�p<�(  � я�DYFfHSdM\.,�j�3c4��>��XĐIN���7�j�� ��-�G:�i>9\�]��8C_#*�v2m��>�]���3!e�ӳ��zX(����%^H��#6��B(���_&=P����~�>�����%�G��7D3���.�=6����&�%�{h	x<�������}�����V-��M],�����m�����)H��z+ڣ�}`��Rv��!��[���>՞5C���ԥmp�v�i-Wl�?�����zٷd��LX�s���ަkj���
>�������{���9��:�_K����iXXt����C���!��W���-�EE��S���1�!y�q2���qݔ�T���Lyh�Z1�i�d�6N~�qu��1'�9��_Gn. f7��c�N�MiI�	�;8:�v~4g��7%�Ye��4IZh)
�	�ܨ���e"��f9/��������%�p���ٱ�h=]���������~�m��[JEp�̻�~jŀ����DKI�9Tt�.�������F������:�j�f�T O����/��4�T���q��@�;F��-%B�kڙ�65h_�뼢Uf�^=ߑ��:��t�t�)Yʳ_�:1���p��ioF-[���Sj�;����go]�@灾o7���z�Ҫ�R� Y���x��:���y����I<9�S��ږ'eN>�9�6M`0�!{�{��2�ì�]�����|.��:�ܽmz��22uWYN�^=m���>��l�Hʟ��v��r��j0"��2����r��������z;ut��b��0.\���Db�������g8��� f>2�h�i����Dz��>p騹nh��-)��:��4:`r��K7?��efD�?����4>~��gy���i��u���``��e����Y�e�����������S�rb��j��Vs�U�"�t3|%io�-� ���[,��[����Ll]p��sZV)[y���٩��r ��lҳ����c�٦����Ww��kv���1���j?�U��F'�����}�
.<2E���P�Z�yM��A�ORX9�|�o�Hz[�ek�Zl�ّ�b�=�nU�ϱr�����T�� ��[��a���Y�z��;K
S|1�3�p��'p��{2���.D���QmF+vZu�!|Q�5�Z7S���U���,I߸����F9ا8���&�?�^�^��<�k=>g2c�K��7ie����d|�5-��)�`�~K�h7��ZѮ�|�f�\*����X,愓u�-(�D#�D�jۺ�4-&K\&�b-�� ��� ���O��Ľ�EE$�0��H:ݗ�i���Чm n"��F��Fr�;��U�%�PaZA�CS�b5EU���5���r���v�,�g��0'��}Sl�&N�`#1�:�.����-���"��Fho�u���K���橂��eh^��Y���<��SVT��5��fv������nÆ�o�&W��uFm~m#g���8�18F�s��qY���$nT�&�B����� 5��$Y��a�.���@��6����r���]}7�g�5u���T�gV�m�C���F�|�4�U�mJ� �����-Ah��$��i���>���g�ɧ�	�{����"�u���v6����x�QW��[��C[���΋L�8�إ/9C> ���z+��o���a��&�U��G�*�w��>Ȣ��n��dFEzT����T ����=��r
��V/C	�3��W��Y��m�.���5�Y?蘭u��f��F3�hD~�~`$*��L:C�D׬�6V��M�;������D�j_��L��é+�l�Y9g��MN;b������h�
�T�.�JO���� #!��˺��F�D�9�#ҝ���[��˻\t���==�������k��!o[�&����5,ؚ��[c&�"UR��>���� ۰o)#V#��C�p"�v�;1���<W��Q`�x�o�i5�̸�d-i9�?������+�U��Q)���|s�N�H��5���)N�P݇QV�3�(L��"���[G,�哬��'�X�Z�G����������2���@>�%�����+����z���T+/��j��&�+�&u����z�U,E��s�H����m�Ԙ����CU��v�+d�V����mS˘��a_�m1��k6������ga|�����MO��K�@`�]�7[�����F�+D�p�M��6����O��.��?#U��T��K��s+_A ��P�)�`_A -g�?'�׭[�nt���;}Q,p�� m���]5��H^R�Mr���@W�k�ZT����� ��D�X�k�q�TҢ��>wL�;�����NЋf�5��)5αp5=5 �D�fpBe��!�c?lN`�N2Nl���t�1�
�,e�}�u=���V�c��lo-Tx���r`�O�	�0��e�� M�v��tu�Ҵ����ڣ�K�޻,Q��&�K-\��NG��i�C_<�	����o���h���v0|\�c#�V˙^���lՁ�������=��U��vb�+?V�9߯��.3gs�,=s�ˋ�PSM��4x��\A�]�e�%:� �"c�>��%�H�w���@&�d̛?%P<�߳j"!��G3f>S}Z��'��B����f~�]-��-��g:ao��lv��WYk1߬t2dz�,�ї�QL�1p}s?�IR�}�CrT�w�v�Q63���0y��[�H��*�>�d��f�F$�[1C.�,��}���;���U1>6Y�<C�)�&|���������zߔ�vH��c�o��'�K���I�L4z�ue�@U(�y��ç�~��Ĳ��U6+��ݦ�c\k�9-�myF5��ՎΝ7���P<�[��R�Cs|߫���>Ƀ��jA��������n�Q1٪�����(|��A�=�M�a��O�j�|\&�G{.Y������y�j��H��:�>׺� cf9 ��k�����eV	�9��cT�3>�j�f���/P�PɄ�+����R��ɲ�V��ܵk�QL��c�q��}���b��LE	� �n�����}����+�����W�,�.ZEd��N��E�Ql�͖_�^o�RR�iwc��*�d�V<=�ڙ�DF���x�4��;	ʹ`[7fj��sc�(�g�E_ep3�a�7L��ݭ����;%e~̵@����D'K��nݷ��r(߽l��ξW1��q��D��O�����x0�S���,�h^R�Gm���م�wm����'?��ۑ�$��?�y�U+�|�+U���]�����Y���0�����)�-P6љg��0iu�R�� �-+Kq��c1�b���?�-xڲ��ڣ�)����vGJvB/l�M��&��m�r�RO��4�U̹����X��T�G�������W?x�������ys�ғ�"��qF�������&����U���[�:����(p���ڏ�yI7��v.<H�h�j�E�oj���mD�-��&B%�":��u�!az.Up�QS��d��F��t]�a�H�����+2T�_�l�b��p�DSPP�>��Z�e�F���p����[�v��5}y��b�#�|-�C��E��qb{-���F��g��i�e��z��c.*���t߫�`D��B.==������+��w,�VWrC�w���/�H��P9LJ�����kEo�_�Y�|)��ST�a��e��	U��NG���+�}uI��:�2�c����!���9��W��̥�BA{��>x 5_���	Y��@�����F���{��V�Hi�o���S盭��mgS_���&��"-&�B��'�u,�:�p�LqOQ�������8�*Gb�����T��g>)�[�Ʒ��{$G��	�~���Rc�Zu���5q�%�lu�Ƈ�q�U˴cD-¤ـ_"�ק(_2�q�9{m�?S�zp`�5=?�|�Km���[��[:{j[I���ϯ�Hcw"E��a ǈ���5���1��W���Ubm`�^K�c�=%i���"�����a6o���|���7�m�/ZME��������U���M2��*)�fA�;SH�C7�BÖs�Vty��N�r����E #�B(�٧����O�����2a�K�`��l���� ��?� L-�G`O2Z}�G��4V�I��f�p�&Ww��ں�<kA9^Q��Wg�O�2��15|m>�A ���@����������QW���]
G�zO�UT,M48�ݘ��A�\�&���*���~>�8�������9��Տ6Ro�RT��T���H�zx�qrr���P��[M�����v:�-:ЉbrԲ!��s�)��{�	F�#L��^��锣2�6�\?�xff�U�D���#��E��r\�|R`���A�a�p��+a���P{{5+��Ic�5Z/��^�����*�rGP|6��t(e!S�����ӮbyNh	��64i����6ЋFA�����B}�b���(�{�y
��<M>���ۈ�
�]]%(/̦0J�f�A~���a��ɶ��rr�b�����~��0��(��4p���	�	\ظ�C��}�{���q�>�˴���mG�p |�Z�#����k���u�L �,Xmc�|q��u�
k�V"�i�bqdo/b�Sc@?aT�#[".(4x��l�sj�Բ�+�u��F�!���Yx6���<���}�5U~!l!� �ԫ���͇�{��	�l���;��ϩn�(���S��������D���-����IZ�f4s#�'�;#��\�ǘ��|FJ{��3�]m����{G���i����/q���3Q1���q"ս������yl6��If.��A�y7�'�)hi-���$�7 f:��P���
�*��V���f��xL��f��0^��+�ݪ�~�^5��T�p'Ł����SfOQ??�`6�.��O]*n �0soq��V&:ﺸ�n��`���Ѳ�-���g��ʱ���k�z2)y/A4/W�wvpk<��e� �J0��E�-��Yg�d��|� �ۃم�����ĀE�`؜6�Й6�xN�	^�!s9>�+ݒ.�`7~�B��MEhC�<2��>����FT!�ʭ���)�(��%x�i����kc�����e�����OA+-طr�pu曖b�#P0�
�hhK�ݘ� J�1R�Ԇ`��zr派FW�ޫ' Xx��f�g|t�����֗ɪ(I������nu@gj��}Z�2�p�U�9%�9uQ۔�| ��S�ͦೇ��q.�~.����ic�}~U�c,������;gj�8��g���lSþ>:�Ŋ�x-�':1ӽk�?����ֽ������MH�!�ZT���,�U�_��i���P��k��~�ey��Vjpvvv�Ϊ:׾/��K8��k8CecM�P���ä����o���bt�b3�9�H��<1�M��u$��0F}�e����W@�5�w�j~|��}H���w�D���+	��6!���/���Um���:�o78�.2_����QM��{��M(qhntZqn��&��r
�(��$����\-R�y���h#2h���P�qx�8����KgCq��*jY��x�բY�����]]���hA���v@v&컩`,9����v[|TI�F.Tc�J7b��:����������H�v����h��b��k�:�B��St��S��`���b�U-�}�*���K�t�Ltrx=�@��.r�I���֔U,yo�Sz|Lz��f�k#���>)������2w9~�L+�K
J.��e3��f�٭���"NV����ySS҆:]���`�ʀ�V;=�}���B���-�w:kNB�����#*�t��I
4/U.�����9ZѼg�*`4h�%����4�X�.���p���"��c�8E���+7ڄ�zbY���@&�G@c�W^�%���$�R�5� Cg7u���&%ëp���,��9ˡ�Y��*7;h6���PJ�}��C\u���&x>�4��s��� ���"�I�Yl��%�6*��r�K\kMt�U'T��
|&3'g��5p��R̡.��|�fKxd���Ϟk���ħ�S&�5˚����w?O��_CD�8�9���L�xۛ<Y¸MGx�.�|���i�-�9=���)JQ��\�5��m�W㹐����Y_�B��Ū~��tb��X� �]c7�X؉+ȧ�� %l=����:���UJ�2�A���c�u������Y�hV.txv[8Sܺ9u�����m�B�S2W��F74u��;?ٟ7��>�k|�K_c0H�E���tW���Ǘ�=Gˊ�X���t
���1`� ~���������e`nԜuþ㑟�C���`�A�M�:�H�xt}6�����yb�>''U�r������n���aWF$�b#/�W��,8�ݗEĖ^��ac�48�iEf�L�4f��-��|�UA���� 3)}��|�?����1q�� 6ɥ�m񜞩���z�c�@rǗ�R��e��2��d��.!�l�ɪB��(|�}vUhY�[�|QHu���0�UHl�)<X5D1�P�m=TR��>���L}�B��|��܌��U����4�^�q+*�tr%�/'W�[r��I��n�D[ ����A�h���0n7��P���}�c�a1p��j֨/(�/��I�s&@!����Ĭ��*�"19�zP��]i�Ҽ;�n��,�?�*`���}�2�>�bݩ�РK|���׍��?�\�^�bڍI��g at �2�)��5�R.�P�q@���f>�QN.����憯���(
�s���u%���6������0[�+�Ȫ�7`�� 築mO�����9svFd�n���!�i�<�g
�UI��oÀ��W��%��$`^슚�W�i���+�SF��=t�4��VH�5�f�?,�ll6�]����5B�50r6H�	���P@�����{!eo�v�xwO�wP�ƹ����^b����(���y�2$��)�j�]��}�;`m96��"z@�C)4��	Ne�)]�Y�����c6�>|0=׏�%�$���9|.�w\$�S��=js~t`oV$��|�Ȕ��j���Z螫]�qv�7�bIN�W+��Q�Ǆm������Mʯ�Gd���5������)��+�o1
W�/k���j�x���+��n��T�]�u9R�q{ڀ���H����U���[9��nT�O�@DT @c��|�t@�Z�R����8@���X�&2H��,9�F�G;����9T>��b4�\L�]!�H��ا�4c�\�e��G���� ��'����'T�EFw�U�\��Z_%����*Y�s3�v{��ټ�ഈg��f��6�<	�h��p\n{����8�I�ᘕ�6��� v�|�Mh#1f!�[�W�2e072��ڃ���vz�>���he,Rlпi��'n��~ޱ�1C�pC�4 ��Hz�!�Ԧ�:�_J^ 6f<��z�?�@ڍ`���߿�]�`��:���iN�`�������'����[���f���jD�f#��#U�PH�Q��0�Ϳ�5m�FB fh�)�
��j�4Q�3�;	�E�������P��Q1G~$���x�3^掟����n�6l�	YU��N�THH�8�{��2�N�'�
�R��a�����3����-�(!�j��n�� ��m�/����r{��I�N��.PC;wr0�8 SLe�I�g;� �@x,)�5 6�U!�������&(��Egu�r�e��Ũ���⁺���@���qmgWAI\]HY]�R�*JΉ������1�	�h��]DCۆ��G`���ԇ�Z��^(��׀z�ҷ�k` [Z�����
@�za+�^��2E��?�@�Es�������'y�"�h���M��2ũs��{�� Ћ��� �Rˢ�H�W�눂�>T�'���FO��p�U��',̪�N���߄�i�g�Us�JKY��Ǧ�ݼ�eB������D��!* 8Ȥ�i9y��/9�%e>r�	�O��{w��p�{0����)C]
+/X��m&�y��d���~��Py������H�nE/bMAkfk������Q��&�6�G@�?�HD���ч�o�x��y�m!p�p冚��k��j΁']B�X�0k�?o�miS���y�v�^Qa��#)N,�錍,W�(V�m�����o��(7�FײY�Y�ذ{���>���Y����h:�����v̡�<VD��>�`2)�Z5ߓ����2	f0yU��7���C�č�n�s&�{G�eJ�'p�OL!�FTf݄��a��ȧ}�A�G����ܨ6PQ��,�⾱H+��%\�h�a	`�Mq����G��`��@�=:���G�ps}+%�䠄�������<E���<�2��e�,���:���,���(�[��(�?o_Ϥ�%J -pD�>�h�0W���7�l��JBe�����v���kT�a��m7�ϒ�1�D�����۬��U_�B����U%qa������4tf),l�ȿ}�S�NU�¹P{��/?!S�)Ԋ�:lOR��)[^=0�+�-O�t8���2��o�_�&3l릛���O����L ������+��BP��5J��&,51�ObH��U�B>-�4�al>����ΠM���e��ZC6� A*,x�|�q��׀��l917:�B�ITDD�)�����?!w�O�^-2����̣���O4�W��b`s0V�REC~6l<�E�?מ�w hރi��2ϑ�jk�PJ�+2(���(�ȅ'[�}^o�ذ6�QZ5�0v}�!��6�u�4m���z�������S��c�� �x��bGI��uQ�����,cas��c���M�#�Y*ڎ�H�V^����_Qbn�e��+S���1���q(ć����Ȃ�PN	7�1��㸮+x��b��<������ύbzk��\���UXq��xJa�X��Y��YGg�0���L7�҆��U�������t��`Ø��b"�Kq��+LćQ�[*�0Q�����>��0P��f��HK �w|�c`C�A���~�ɣ�z&�����l���Ap}���Ղ	�Mei��?\��4|�d�Ūry�}�RcI�w�k����1$K��PAcy����� ���7��ø}�xT���#,�Cn{�I�Aʥ�v��#�D�1�!�����^*%���?�ry�^��!��G�!����t<��W���}Ǌ���oU�}��G�{��G�{��G�{��G��z���d�*i>s���pw<v�髧�\x�j��������[�y�ݻnO�M�����alD���y�$�K7o_?y����'����@<:s��Ԧ�5fĂw���Ժ.�o����C��w~��ߑ��uj�'�w��s�������\���w����o�u�_��u�_��u�_��?����ƪP;��gu����Z���@Wn�󪴅���2�u�ex(��p���H��?m��������Pΰt���m�A�){T����i��7<��a�M��*7�V�)�5��}�>��ψef[kI3n�P';��sb�����vͰ��6�"r����&ް�4'Ҹ�E�ӎ�w�B��9;�Ny�ï���@�X�|�=7M�Vk��aA�����.޿�
e�)���F�{��Y�Y�+����X�Y{����s�߆��i�%�&Fx�0� ƎW��X��\Tl�p/]�m�Ƴ,V�q>��R[)g��a��REգV��n�L>-BU�b]�4C�״j�y�F�<i8:p_�I����-p+ݒ��*vCgY�8;��U�;,������&�r�ѬQ����Z��ɠlPs��J�.+�W�uKz�j󐹺񘲗	a�����d&?���[�r�}秌Dk�:/�!S�O��6�_`|V�vS�����-�ԥ_��#y��!�KF�U�H4��,�D��.��<�ʸ�E���௖�1:C��"�������_�ɺ!�Q{�(vZM�c�?�E�Q�Q�)�Pc_�~@ƌ�UƠ�^��n~��D�����a��O�2���Y 	��ӈl��Q��hR������_a%���0Q#k��,��e���W��sC����"������ +>ѓ���ܪz�Y7oų���j#E؟�K~��g{mk������	�79��n0�[/����ޣ�úE�G��-V�D�D�W+��jQ)���������)ۮ����Ȁ�]{�7�%>��ƵVw=�hr���2)��;G�$�	�X�	;>%f�m���18��2L���}���6y�W�8ԥ��Pt���UPx��0�w�x��5uGч�r��#ĳ����`����rm��L���:��v@H�I9�Y��:^�s����vU'��:S���i	8�bI��S���ִ�zLo�f��L��Z�/�{����^��}�jc�{�ʚ}�������)���l���⮎B ����y����qb�8�������S��b	x|ӞƇ8kIci�Z쇲��8�S��x�ύ�VG�(wO�L���5���:n��?̧
�oh�m�^��fݶ@��t`3�R�-���*�#�kKӱUS��jf�j��6G��B���Bz�I;<��[����&�ѐ�b�R���B��/Al��CT3��}��:KT�x�ۡ���,����,�C�)sGN>!:߶��s�_咊����\o82`8�:m7L���G�����`�g��_���ߋ�Vq����(�af�ZE�U���پ��,��o�e��xz_S���/�x�����8,��Yv�ywuY�K�\���aR@��h�Ӛ��Uk��xņ[������m���{U��S���r0�8ê�H1�Zշ�AzF�U�������L!�Qsr2W]\P��k�\����k�v��rC\B�q.�ߊƈcV�d}áS�kg<ZA<9ΫuO~��kL�����c�3�(��̖�`��n蕋`7��A�.���쨰������4L�b�}���I������c��Ɛ䔖�5�5�d<
#*Vo��?�����cV�O�mG7��̵��"���x���ъ #��5rl�&2��ͨ�ql�_�<�ԏ-t;#|4<y7 �b�M�|����B�p��S�lW�+��
���U�,��X�w����[��Q��0��S��p�OԸ��t�${T���_�~�,��Ʃ��	��JJk�N���ʶ��TB�ZT������@�`8ꪨֲ䵓;�D..��_�Ihm�q��괺���`�����½~������L!�)�@��(E���A!�����k�l�R�qGL��e�:.2T�v☸7�}�#���E������9)��L2;�,b�~��X�-p'�7>�Go�JnĆ>�W^ZLf��#r���^*}�0��g�ൗ�"ꚮf��w��
�R��[]�5��r��}��	����ު�"8��`\݅��4MM�C���]�.�R#E��� >�a�<�8uJ��h��0�yQ��[��ni��JQ+����e�R+{�f]�;�#y�'�+��*��I�>���p��nߣy`��M}'�\D�*cp�ӦSd���HFd����Ŋ!z%7��|�с�P��M�C/�%q��.N�g�CyMuf��D����poh�U�������(��:㌈����ݝ��n,:���gl7�����P`$L����9k衙M	�hu��Y�*^-i7�I�(�`ts�.%�I�^��^ˬ,�T����ՁoS� =����z߭��?&��m��;T0���ww���� ,�gGI����̾�o�ޗnx���bJI�g
�LH� � {Ă�B�r����,���%\,,%���ػ�ܵ}g�Rjt�*â���@�T��ׅM&_���L���׽��64%�ؑ쏽>��y/�q_��cS���6KO��U|lNN9[p�t�qqysRd�@Y��`���}��W%w�1�U[h�I<;QL�zsF��[d����3��l�[5��o{($,�z�	���:�������3*�E�0���4)!:�  ��U�� @PFGMZ��J���C�C�B	Bh��s��{뭷�z�}�}�bԹ7瞳�޿�������-�)���a����]Bs3Q�=q»�n[_�1�a�u�Ij���.o���'�=�eN�q��\�B	�Y� �a:V��$�ߦj_>H�dX#�Yu-��0��u^]Ĵb���ri(̤f��UÙ�ϵ����gS�jN@_�{pyV�˴׳�os(��7�x������97U�	c�-�{$�R�tpآT{�u���Ơ��#�Zu�A���i)؟�+�k����,=2���G�Q����@7Ҳ���EF©�SҰJ+d_���dz$���"g���k!~����p� M���+xS�h�s׃�h��@��9���h�'%�Wf5;$:�cQ�����gϧf7A��vH��̈MC�X���f�g ��+am�ۘK1
�=�e�������k )�f5ϖR�ʕѲjy�@�@��Op�����q��<�)1�;)��k)�˂��w֋�@�^t߸��S��2���c�p�i$�4l+��;�w(C�g:��NO5�(��uR��q�	�>���A��A�~���=�T��cqi�'o����F7������.({�mwL�q�ˋ��'�����,�B��G&��/&[���5y�����Mz��Ӂ�Ʌ}��v�e����}��S�q�����h�n"�g��D���&��U/u��e��*��h�d����>٩A�&��M<�UP7}�z<U����<Gxe�~�V��sq�6뇄~�����/��G��4��>��b�,t�t�z��S:�1�9G���X����A��<�o ���(����x�wj]��»�Tha�Zm�P������A�Ó���]k��+fR�*鵡# FmU��|�@.�ǋ]LN;���}��+�OT�!�)Ǿ�<-:ȉvIe>������Kx?9���!衪�����VRk�*z�Bh�h�h]ߍ��4���N��%�D�Y���:4�8/�UY0K�sUr&�˛7B+7Dxp�Y�ߢ��	�._z��|W03�2�=?{���l��SST>l+���o�)�lF%�*�0������N#_��	�Bw̣�J�]��Ns`��%��,�$��������+Cv��<`��_��Ռe���	 YU!h����S���.�f9Kj�tb�3^��~�]���ǔ��yWDja>G[^l�j�i�^.�r6e��Vu�ʧk� 2'�D�����b�Itq�p������?�^T��Gͼ%�K�����ٿ�I�5jW��w�\Ŧv��"
nǵ�#í��H���Ͼ�H5��*����`'�,y��2R��o䢴lo��%�Z�]�.'��~���nk��P)ۈh���<'
�����	x��ϼ<a>k#[h� �Y�`�w:ђ�z1�q�������U2��eV�z3Mf=U�4֗$Ux�&Aq�/���t�k;�
_�4G���l�9����"��֕q�%��Nk%9�L湉��fȩ���\<��Һ�r�a$S���*�"Q��-�&P�|�O�(7��p��x|���>���C�;�t�S�Z�f��S��ڡI���T�����򢧺z,=z�����]=�\j��'Px$��ͥ3�:c���*�d2����k���뱫�������١��kG��oXqC���^:�X�:�3N�Ժp�ci�wn6����[�'���=Pxib]�Z��	��_͓�g+�*llM�w�h��eq��_�-�+[�5"T�Q�W��j��p/M��4� �w���~��$�3�q<\<��f��L�ZHomp��(M�t{���:6;;�c�p����e��ZY \'��M��&1:��{�����3��==��i{`B�Y�R���w��$�R���A�=G�j��7�&�$�k��n<ʪѬ�s�sï<.�%M�X8VƳ~^�|D6�2\!�S-�q�0�L�s2>>���s���%B�}��\mYX=�Kԟ�y`,��?����qe�����o�=�
���{jn2#�B+�zC�!5��k��ķ�	p-X�|����<�pe6n/�F�~z�ǎ��f�z��E�GSav��i�c?���9\�l�]����*�A�B���q����'�mݥa��U2M��H��I㉛����1�e�Z�'+A��rx)e�^�MzvU���D�z|�ΗT�����-��f����V��.�L��_*|�H������&�f�A?t~H�.���|/�եs�4b�R�6�"��ٳ�:�.���n*AM�����	���f�x�Il��Bz0��c��\4q�B{�RC,�+��¶�ۢKz�v�Y6"���σ�i`��������l��|9X�mq��,��I�2%r���ښ�(�1'2%�r�|��8,��)a��t�d�&[�Ǒ
�煛	�Zu\�o���4��x����އ�k�,��v��0�
�l��Z�Q������i����AՂ���xT�Ǭ�9lY�IIWᙀ<�"�y���8W�����R<$R�H����u�y�����là��Azk�f�	n�L"۵�����6?,�+B.�5��!�	�ҧ�8��ۥ.l�����yw�Ⱥ����ے��C��#�2���Ƭ�M���AhLN_����MaINx�2-)��y�5�ϫ���&��=/g���J�H�L)�e��+ �f-G��2l����J��M\4vFe�Os�/�7m)ּ��M��@eE�d���^�H\��\ZZ2\>� B�H���UWx�䀈y��}�O�M�Ѝ�#�B��g���&��!�9v�ֱү$�Ѱ�3��F��:�To +
=����j��74,\�z;E�$C?JjzDq4�v�A�{$�^������p����4CGML�톓��� ]g�KZ�F��CQSJQ�����
՗�S���<UF��p�U+Kr5��ۙ�4�
�nXܠ@���F��MK����<ԥ:/ٽ��
3Y��P!FĲ/E�y�S{���ȥw�V��o�e�	F�J4#�K����&0X7ڔɝ?+��EYm�OBx"0���h2�<\��Q��#+c�̓�=�� ��*k�:��oJ1]jK�{΅����N';ȥX��xű�!b0k��I[6Z�8݌���c%(p3r�"W�Y&��!c@���q�,D7��<�)Y;���O����܁�[�x1�VD����������@��TM���܇�%Av�zZx�a]�H��M��-�g`��Q*��.J53�|V��&���eEfaWt+�N>:�T<C9P�!0�A��ۓ�Y����!��Kɭx��� ���+�%O�+�Z�͠�`�L�,��K���5��e�J���<��6�z�f�����E�[0�2hǇ��=g�J�C���m����������y-|I�a������գ�F���F�Z��^M�k�_-����2^<�^Nab�i�-D���'�����\C~7�fO�+S*��.�x�=�R�p�8�`�a�;���[�ڢ��!�؛R�H�E}��H��%:�҆���"» �� �_7m���������5���	�k���F~�f���n�S㌬i�/��!��^�x�N�,_dII�V/�32��e�����t��yݬ�s �u'u�Teq cH�.�iH�y�_=����H��m�H��U�'4{42=fّ��k�x�Z��L�X�!L�)&/&I�F�B>5k�]l8ue0k`D@�q!5��b�����V��r7��%�{*�f�cc���}��9���%�}{i�I� �X߶*��"
��UI1�ި�u?����Y�g�E��
g�Ck���2�U
�A/k�Ҥ�dk�t)�i�oQ��dG�C�h�c�ZF��%��,���7�C>N�ΐ����)��s`B�0S���^?|Aѽ�o�٥��9�	�h��V"K��0�bD����m�ft�!9q�$�9Ѐ눠��xO�����Z�ݭW9�젮|2�=-�^��W=�[�`\�m`S�����K��d�C�j�/L2����J�v�5�ma�9�_Eyϒ�Z !qkdBt�"�ب��y�&`�`b��*6~ձ��Yܰ�}k��2��W{�rE6��?�)�j�|667����`Z0>��v�yy�P��^-KV� �*!
�̽K��qb0��������G��tP`���GDn7ν�
���l*y�����ّ�5�i~�ٲf���4HP����&B=�i�V��Ũ`j��=q�-57�w�b�x�Ih��+�!�At�|�{��&�$���Ւa�6'�4V�������||��롞=<Iި�].
��@��U�0�0ʐXD�nfg�]s�I��>��,�<݇���p��$��8�P��K&8]s��ރk]#4P�p��r���(�bj8��_�����$+/�L���,y��om��t6Z,8��B�W���~�8�����{(O=]�|{��j�j?�����ٷ:��"Xk���p�y���҉�Z��̡�O)\>���q�k�0Pr
@���*�M�6.�w�ef\o���5/9��%�B��$]�I��rSز0���zm�,�n��� 롍�լ�li��\ ��ǖ�-=����h��fσ�l�j��}{��:z�6}`c��m놁����Et3JF}1+��j0獁�q���\
������$FF=e�-�uH��aA5���؏�J[=G{.��1s�L�2*A��rn�YV	)k����ò�}�%������S�n�H�΀���0��ᗻ=4HB�L�XYV���8��T��V�e$�FB�W��҄��Z*�}��{�6Ҙ�k�(�Vq���p�^Z��O�ƭ�/�%�0A��z�P�XSB,vU���~n�I��y�}�\�YiJWц�\����?gn�'e�j�s_�����^. �vÄ���r.|ju��?��yiY����C4�L�iM�o�5 ����}-w��9͌'�C�r�����(c~T�|a�����4�ݰ�V�>�a+��@�l��S��S`�!
��0��%�X��%�_��R��?���S#3�1�=�v0��؍m17�G-�����ا	|���� �0��������
���l��νUAg��(	�6�@l6o� �#�?r��m@��p�S�����1';VH4�`i҈�҈
�|����?yL�l�zJ�'-J8iC�Z���[+����6|�m��X/�rڭ��t����Y��ߝ�V��}s0SY�f~Tg��	�P,��������)�f��(��J{k����;��7G�M&5^^��,ڰ\�!�1��oA�&Ί��*1�xh(�_\�u�T~hRc 0k�;j��ve.�2l��vi�]q�}J�)(n�jfi��z�"�2 �f����d�P�\Kߵ��@M���1tpk�̣�y��]|�c��Ex�����`7�1��i��֧�Æ�P�V	cAˊ����Ez�uHK��P�{iq`��䍆Ҡ�����۞�FȐ���0HL�|�f��ۏ�6
�� �4L��-�m�]�'u�&+���`;mh��˓�)=R~-�"�;(U�գ��2�zՠ�/�]s��1y���͇��;!2�W_.|�z�z��<�ㅣz ���;�h�i?������%�tp mJ�RP)��C�Qݧg>���\�aU(ϱNW�b�4���m�2��pVm2"�u�Vm�X�z�U�j��5��;��)��.���	����S
��;/�JBO���WDjF�}�2�*I�o�p���:c�#5OB)Sj|�*�L�9����Tc3���{#������3�Sԓ]��`.f:*RG҄�<�8S3��myDnV�1�ߑ"�Ir��523����0�?aH�6�X�U+D��d�8��?x܀��Ɍ��g[)���}ƶt��h�������:����m˧�\���}�jt��w�z�5����Yy�fi��{V�)py��m�ʮՏ��
��4�]I���RJݙ�n��Px&�6FE�w����g	=!J(7����Gv����jz��C^�ʆF�3� p��|k�|�j��.t	�'S��+��F�-��G�j^�΅ջ���%K)�%7�w�y��J��C��2�t/�q�=;�b�wS����ڏ�)6�˱��_�{��"��8�����ӭ��ӝ�:z��Z���K�/��{w]�~�|q7>�㎨ݰ����#�x���:s=� ��$^zJǞ���@�/�x��mm����A���5� ��"�����\��b
%?��cb���X`n��L�f�ĳ�Xi<F�.<�ۮ��t߭{X�O8��f���2`}'�C|��K�s�I�Uσ*Y%�:�%�×F=8@���I�`��Pw݅_ݸ��Y
3�,_ 
Jo̔ͅ7���G��hWв�r��e��j���F� ;a�2���M��|.���O`�_9D��9 ͗�:&��&$5"e��bG�]�t^��ruu�%7�����/9b��#.�������
Ƶ��~�v�X����3��y��w�A�����N�m5�ӕ��#Naɸ
�������ifB1��Q��;���,J�MH;"m^��r��1]���t��Am�Lw��p�i	�γ��+���p�T�P �)Q��ݨ�����C�ye�.�{��=�F��@�GQ��ԥ֨�_���5�G�ov1<�U����E��-Xj���5U���-��Ε�K��8Bv!T�ܶ�E-"	��\��hU>�T6OO8�ܦ�k}��θ��v�0���.�b��UU����gO0kR.��V���i$�'�ð̊�UF��'{_���>X�F0#��L�=mu��&��v<9g<)qYbTY���l��Y�Ǣ#Ӆ�!6����]�A��D�����Q�IM/a��չ��vž��w�V%6��	�=���"�P)Ê�9��Q��Ln�s�v��j�fx?�2A��6�J;�Eb4\k���4M8�р�pPO�N��q�[sR&դ�s������&D��jE]zf��y��#������}a-|��I�R��RA;t�/�9�j���]��Id�'����Ȉ�n�4���m���c�KQ1�G�ҙ|M�*������A]ݞ~������Ƀ�b&�.��h�=P�J�pԨ2�'%5��.G>����I(`��O�g#E��+q�۽u���n���u���U�r�I����s[}=��G�����L�*�3������N+���`����3mMRJ�7[����2lF�l!U�x���~dF�H�K����kVf
�͎񷫈��x�c��2ZQj��B�ե&X�':8L��T0%~~<�"b��Z`�ZPf�z�������58��uY�_�����ܮm{A1J mH��67[��
�\��I;q��@�è�S(��d�#� � Δ��p0��dU��wXDB-}F�a�K�hK�▪'HrA5��;ov�����=�M��h�!Iv^2f,l��ԓ��jX���hA0��*8�2��5�c��#sd&���̜.�ٿ
��WV�+$r�y�see��0P��h����R�i�{��}<N7�Z���&���F(�I#ώ��ڃ�nMާ�lk��/_:�ɇ�5P���3�Y
fɘ:"҂Y�͜x�F��A{y��$Vu��%�y�L[j�lA�x����:m�{�D7�P���	�F������sI�Ќ3��@S!���'7Y�����w��V��bLF(��Ӥǧ+��q�y�ߝ�y��̐tyRԋng��1���v�S+�&h��4z��
���D%S�s�x��R��m C�����9��pc,�<����O��	<������倱�⢀����r��G���+�ِ/u&�*�;f�,��#�e�Mm������i�Z� B�$�|������2*?�9�LX�I�>�#|�yMݼ���C�*k��o�D:q��\<Li0cqD�)��@����^�:Τ�v}�b�*��F��u�,�f��F�U���&3��"Q�J�l�3�A��p�jx�ج���D����͊v�5\���Z��� (�HiKg84���x��u�U�3y���%�Q���O��x���b��o{-=;���6�W1����\��5���s�S��\Z���l9KF�$�u!�V�TV��$��M{�E�)J���J	�M$/7[�T��&Mg2V�#7v�g� ��d�B��!��������lB���~6F�o��*���d���ע��`�Q����1a�78�3�*E���{���ZI����[c}�}��;�Y��ڦ1����2�'���?!;3���,�z��[�mKfJ�����G/��4�x�9�n����&��p�˼��o�{�F���&���0��=6�%�M��/���*ÕŨC�Ze��!�����L�-p��)�Z*P�iWt*s�G�P&T�b��ez��Pb=R]]���W����г�!��p"�J^-O��V�$������L��e�?��y��e�q؆�Z��1ǥ	N%O�(ti��k�ϝ�?ˈ�Hz�v��y���iu��l�'��2�ߔ�n����J�>R�����4z5�6G�e�Õ�Z8J�X��w�A�\7��INS�\��ا��e'9�?�Ӳy��^�os�fu3X���a�'��C7�ˁq�������s/q�V;��J��Fʫ����-eȹ @�.^ץ�Ƅu�[�"Tu��:�5�W�:�Pm>����u}�o��z�e��G���������ݞ�4�\wrң��/�Ϻ��<����n���H��{�/�������C��"��WI��yz�	�͍1�Q:Oqn�a��EׅͧG
<�����t��̭�(�]�j��Qͦ�YG�/,�>f(�C|�in�E~A��ݼ��/H����d�5��Pt���;�¦��o,̬�W�>�6�*>�����C@N�(5�P9��=�3������]�HKFʊ�Tl0� G޴|Ð��o���;ب����3X��_��nQy>�aU�q��nG19�. �Uˣ�P����:�C��[{yH4M���"'�?B>�B�N�1��2��Tu޼N��:t0Y(h(=n�o�4|e!\��E�2���U�W�w�?�f~��I�n��'���ouW=<<d�-�t��z�9��K�$P8�r4���P��N�j�����X2�]Cx ��<�|��˽���%z�qC�j�A�{Z/�;�MUF�6��1��[Ve��e&��&fK!��u��gn�?�|�Vfb�;�%3�����$?g��2N�XO7_"5�
�Y�����#W������]��jřWl{Ff�����I�G�����s�E�+��(��g��V�)>��"�e����[��Z�1w��E|~�REP�wk5Ŏ�T�)�2��?���\,У��pk�!Y��?̎�|���i�%�8��H2�ZV���ryb�b�*�a6a�3(�}�ĝ�_�0����O�e	̶?%�� з;#�e�Ƿ���+�} ��S�P'�����v˶��-�bh�����j��.묚HLr�@��;,#~�X����Yr)X������$'�ܬ���%�0�U�J��	2�V[	�0%o�Xe��/�ěz��?hxb���b*D'UB{�\����T��B5�����e�`Sٮ5s|RM��z�y㼋��[��B@Wϙq+)�	�,��t>���N�QFi��uF6���P�=-��-݃�;�D�K�$T&8DWu�1�鞝������_f�ХPB���|����Ͻ'YR�j��35-���& ��f�������Jc"��S��ɏ����yz�Âǎ?�FBI��k/����f�~�S�CM���h��v�tc@.We�O�{�%�H@�f���^H?첳ݓ��PG�U��-��9K�	ր�"ʐ�?���c�*����r���p4�Wtm{Ո7��V�!�<��ګL�c{Ώ�i��s��]V}��#�s���,.�#c����<�������cew��Ju��~��t����xlkr&���H�<�P��6�.��wq��ᨋ+�m�#S�w��(:ǜ4$|�p��r�L�dwƣ!*k3�̷�p�*��~�S	 �Pm �����I���̩��Ԥ�V�,��kC�w���1���QT{�?��?��i�lh�	���nd
e_�O�y\��|�~f��b��!"C+�M�uM��&��^pj��x��OT]�@W�v'TɃZ��Y[qZ���Q
 ��pDU�8�h@{v}�i� �H-<��͛}"��RP��&�����
� �?���ӝ)r,��!ny̲��{��C-%��(@E�Lo�Sp����w��뺬�jb=L�����b���Ks����vq��[�	?�#_�{Oc�//zI��y��U9�t%�$�DM�賐���M���sRn'W�q�TC:�*�[t��*��_~�=7�˲ӡ�K�3s[���дٰ�ͣ^�?A��O����/�~l��g`�X��īh�y�ҕM�/\���#�_KK+tmHd��Bk� [��*1��fyAF��t���MkA���F�?j�d{���$�F�?
�gJ�%z�;S�1W5�;�>	��O��}gR�m-�I�"�8 aO�R�k�u�4F^��H�G���-�N�=�nZ��<����lb���\�g!�G�_Y+���O�����$(�f�ws&��m�,»~��cNx=>�+��	�{0�3╓�����4A�	�tt�YFF��Y���4�m��Q+�ޓ�2־�#~�k��b�n�oj����
m	�ҾZ|�妣��w��Q-ί"�'����䂄�SV���=�����'��n�a�Z%ه ��bk�C���q��s�'KY�x��� d��	��K5Y���EA���.�aݙ<���І\O�8���z������c��N�pk�M�1X�q��F6���79��[�I���f�|��Ӳ����|�T�ھUm�
�m��ٍ:��8��0���B!Z��gO�x����[��m��O�W������"eswT�k��Sj��A����.���s�l-8m�;���.�i��<L^F�|О]0�i�';-�q��fe��>�Ča�r����$�@>w��O���
���R���v�bvš��q���_L��r��m'����\;��x+ܥQ���%� �	0�}�g��j��,}�Ҏ���"��'�;���G�#�;�����������F��L������bPR��y�ި��ޭ1*4�X�`��.K�}���jJ�9~g({��̢E	m���Z�+LMlgjJ!��PS�0�ב�m�����)?�aǠBω�G|�|�p����&��Đ����YH��k�&�W_'gV�,wuo��&O7��%^j�^�`%F`�������V��݆���^�+C��T
�Bm���7;��?;b����ۻ|�6��H�j��e(����b
qK[���.n�i^� ���{�#�do>1+C)ob�l4�d��NL�I���=rP�*��_��X����塋��%Ոq����P�\�EU5U���K+�n����3g�&�I��ѭ��Oo����*5�D����R����~�f�χC�kVѤ��")����k<T�����tF��C�8VF�N�|��>���7tv�1���bT��U���Hql; ^���F�G�,SS���Ѿ���{x}�N�tm���|9RqUs�oW��i���Q����2s�&gܰ*��������o�8t\Ov �w�O�Z�������.w\6���{��A���0 �P�; ��7 �k�ĸZW�տ�?�xܿ[�=j��!��_�}B�\N������5
�4�[_hi�)�rX��-����3��0ٛ-c�Q�8Q�CJM�AW�Z��k<�/	�Ѳ3�ZG�����WpJ��pٓ��V��K�?e��Y67�*�W��ϾҪ�9�U!UGD�R
�?w��,�M�rJ9ʙ�T@4Ya��К�W-���q���kֺ�&��b�� ���<��z�j�Ǻ?�S���^�����&�YR�	�����F�*Sj.K�6A�	x��x���{V|:�iu�',#�_��5�썜�Z����8ϐn��P��Bs��|3�5)���g��ɸi�Ni�w#L i"��n�>(G��}�XSD����b0q����E\��X�vRr2�6�1����O�+�ε��o
��tL�O����%zF�"!6���o�����rn����#��i��)_�2���T{�s|ƜM�M�BW�v��m������H)�Z`��L���H�G��Ϗ�nW4=�o�8�;B����SEU�s؏��F��6Uv���;foN�n.~�1�V�>/�|>ĵ�{�����ʜ5G�=�^�Sf���̂���h,r�z�+��8@k�`��̗�LJ�u��c�q6f�2�&l(�5�&���ۥr~�0H���&x$I.6�u���9OǮ��8�6�{	�?*��*�?�T<�"�W����κ�.�R�f}�E�̒����⌦O���s|��/g=����H�Ν���h���l���I2"Xc�t�v�G�32���$��
��/_�ZЋm�y���ў�Vt�������;�ڏ����Ô�`���U�zQ%s�Q�l���IU>6%"(�G=|��!~3����Ys3�M�<Ky����<W���v�i�%ۏL9B鳨�OAGf�G^� 3�i��r��A3�-z<S�h|��_q�n�4�I�8�j�Mni���gK����6x�Ǧ�A�)�����Z�A���e�[a�]�;j9��D�L�ɂ��`�����H5�z���;�=Q��*���,⫞�|Y�M>r?Ī蘤�\�9���9�������I���z�w�^˽������X�Y�Q|1 ��'[[>���jr��D�%�H�&����v'�W��h�SA�F�a�W��[�.M�=�{�8���%/N�SD�Pw_�NY��1�y��T�����lmp���z.R��\��B��3n���|^z�QSM̎y� iȪ�S1Йf��I�S��f�*ڙ��I>4uh ᄌӰ(�ܜf��g1�F9Ү� L��z!�����L����U8Pq�0~���g8���nh���\[HT�q�
\^ZZ�kMQI��C��>ю��٠5u�ؤc$�BQz-���3��L�B�l�Zi�D�pp�QÊCL��q��[ -52���s�:�����l�P�SF��l���0.qq��]��Bt7��9J���9u�-�"�<���\_�~��Р6�D�:7�2�fo�M�(���mE�}�|���B��
tz�~C4��:\>��`�����˜i\CX�=������EՀ�:G0\��7:���4{���"��}��Q�\
B�?l��}ï�RA^�f�^e9�@�$}7ԎReB�##R�f����I�	m(?D�ML�<�;G��ɉwC�z�j��z�Ք��@��{�p#�+vs/�"k�</�VJ�?���.u+34t�;<4`Б����1���/�c���ӵMxae��>��2@�1w�\���K���,�T����&�QFϳ�4�)�&������~��UO-kYe���{�D|��+�qI@پO�x�nߗX�:)����FY�W)�ǆ�*�ńSNhl��9e�xbU&�z����薠YDA�#̿]�$���(�Б3��-s��H����PmN�۝T�P:O���?�F�	�)��b_n��X4�vvj|�|M��ֹ��f�R\��� o�����F�Ȕ�U����	����'l�:�__5��/�VfW>1cRI��Lc����R2�� $�FTUU�ǟh��o�E
�0�\��O�}d1�80���|c���e�K���q����O�r�ci3c��d�p� ����
�B���C_��e�vR�zv<\._z"�UG_*�:0��=�Ԣ��hN(#C��m̂��-O�ҕZⵚ�qi���2�ʼ��U8j?a�������(��Q%࠾��͌yA�l�2J��+^�u���v���ߠBǢܩ�r���&`A�	�*|�_.O{1;r�����	�Nnu�(W�瓯�K����LW� ���(���cL
�����7^\���WWWg�݃2m"�����n`�^���~����ّ�O�u�*�N]]Ă�-����|�E�[v��$Qp.��V`R���I���T�%���j��CY#_ޡ�,z�� ;>[:
�[}�o|��7�h�D=ܶ{�*^�z�p�V���#�Ň���������;����H��Ώu�/�~ �X���mm�~P�!�ڦ��}V�������+�p���2��eLU1؆��������ғ��%�k��g��������wN���t�{=��<��B�����I��:�����W⪁֛�#�H�k)_�8�|��W<;�֥:W��مW�U3u��l�7�`.���HD>j�b��bD�=J����vZ&���5�w�b3�: �~���� 4!�uH�`��N3�Ը��;�7iGz�_�@=d8i�.����X���E~�Xًq�J�r�Z2��rWV@<'o">X=������c��X��h��d�b�m�1��ܵ��?�6R���u�c����5��������z頿�5���vŭi����*��y$����}���Wk�J����O�4�}'WI�E���8w]�^��H�M|���`�X'�X\��aD���*֛y|��I||�B����)Ĭ��j�0�㾜���n�*h��%�T�DY��\tu> ������������.���I=�9����V%�[x	8SjA*@ר��)�$~��%m#k0�Zd��p]ЬZ��D��4[���'��R�H����w
uȒyj\a\�
�Pa�wȳl(S�Z��Ed����ON��Q��G�L�G�n�e]�����Ή
V���m���v��,�p����*QlP�flD%����i���t��x<�\�Ȓ������M>���<3�hϓ�*T%�R��Y�s-p=�sPPA��ls�M���"��'}��S���-��V��������9�	��}���;R�&?�r����1�����k10���[��f����Y�VhZ���qq���Q�(�q���ա��
I����Tg���Q�x(��Qb:iG-��lk�����~�'Q]��r�r�*w���RU����A`nK1���zg{�X����Z_N\�7��AN+�6͟������%��wnJ;n�7�7�����IU:G�I j�w�.����'0!fs]*k!�KD�|&O�I[3��� ����}p�*���s.���).�h�;ũҬ��g�M���t�cu���\d�)�����F0P�p�o` �1��q��N;W̪�wsJ�	�5G�7�+���?>�m����'��.��P����B�J�����]�"ѯ7�H���r�bϞ"�]༂:
"�;�p\���"{�����e�:|w�_y`�������<Zj�"2N8��q+X\w�̗�b;7����Ytu^ @�i1f�S����1�@ �os�۶>"�������b������D����Y&�$ι���3;N��K�[����s��v�H+$L!��Z�S �H�/��5�iN���	�9�h��u�WJ�H�[f�)]=wj��sSX<�/���g8�5�'����#��nc�bI��?N*��`B2uu��}bM��g�j#GdZ&�3����
���+XjI*a���h�~��OdU��Y��Νu}@���ly�� ��0vn��:�T���q�_�OS]�����g�����J����us^T
����?;2��nI��6�ì��y�	�C�گ�}-B�V�<,@7����ů�yS;Jw1뛕�z-UV2
V������LW��V̬��O>�l@u���S������>/mY|��q��(��o��.̎G�l"o�jz�[������@xwG�x��|t��΍�C݅��}t Ɉ	>E���jSՔP9ۄ�:n��U�6��䀠@I��w��E#�ɧ��ړqy�«e�#�iG�qLȭ���m�~1��'^��������1��u$����n�h%�p!�HD�!P�;���_��Ӿ���u���m���xj�
�9��@̰����XtC���5�j^E����q���׿�}�7��03-9�t�����ʾ�NYp�=H���1�q�	�4��{Ay������U�4��= ��y�ix.�e��0��9��z\R��=������(���������*��Ϥk�]#�~*z�������Ύ ���d�H>����i��} ���'v�C}:�O����'�����b�(�2Tv���ǾdQ�qM�=zp��i�����9i�EOb�ۑDk��Q{��#	�^����uk��Pe�7 ;��tHNQ�xQ{(~�D���tc�$�����|�����<����%M���r�&��sv點�$2c��:�M��"IT�"������s���E+%��k�[���JEQb���օ�W3h�5�4��g�qqǠ�Od|t�O�.!.�2�D/}���b�s^���P�K��G�bC�z��jD�o�t�?JW�>�]��N��"��A��� U�?h�+n"�9q�M1䝦#Gn�.���	�U�Ɗ�xFH�Ə('l�/��QO����Z��A�|���m���f�C����`����ŉ'�B�ŵ��L;�~S�f� [䫦t��\}߱�K��W���n�z�8��� #-ٝ�j��\�L�o��'�����%�ݲ�;/��Ɗv�����z!���DE��b-�+|}����?��ۙh7p� !	7!�N��r��Нi
�
.X��
�j�'�jBL���?V</\�{�Y�yZo?��9�� ��Z�?���C��ސ�j�%���s_��Z&�:��E�Q9��&�UO/H��س�fV��͏�w����&m����O~W|���?z���_�ЛJ[�.��������-��Ak��ݪ�k~��]�[��:m��z|��/��o(���~3 ǃ����256�Z-��R�3��a�t:3S���{��ĖH/���w��S���%��~N��A�ü�O�;ֲ��/?u<q෺�����8���u��y<�CM�~T����})t&�Ǻ@Ba��r�bҷ�`BON��]Q��j�_�b�M�M�-���DL���F咤����
�aG���]T]���T~���-_?/�n��p�ߍ.y������◝����D�����^4���}�뾿�뛧�*��E�9�4�3���¯ߍ���5��~�	ɯ����ؗ+�qm�l�ݹv�'�R��3�~f0�t��8�|W���@���/�������;��q�#}�Y~����8��D�.m^�I͒��f<�b�ҳ�/������}K
%���k�Jz]r���b�kЖ�l���vW��́߹p���)��A�����[2��]o��/���������w�[u�G��R,�Wb�֥���-�w�º��20�gN�`�λ _�;�1�������3��{����{�v�ϡ�;�{_e��b���� ���(HH�JKw��0�P�")=�C# ��1 �p��'������]��Z����������>{��+�)g�,����ښ��ɩ��G`*�̱���8��6����������ڝ��Y6l���6���?�Ly��MC�y2��.��|;���C��V���C�n�\�[nш����Q�a�B}:�@��3# I�?.�*����PA"��ѯt=d1�\>�p������V%�S�!mH�^H{"|���T�e�D�e�UT�
D?J������<y���C-�\e8=g���Q��ﶯ~xȐ**i�ȩH;�ˋ�Y�s�eG��ƣ?�	 ��S�Y�<c���I��ڰû0��k<����>D8n����Q��(��_1�.�,4�e�:ҞJ�* �lH�5kxj�p÷�\� �F���~H7\V!O~�0�$$;�\����UT�����9z��X�R߫���7{�����|��ON��7�]���
�Tb_��i8���Η���� z�1B�!��Ƴ�&F�	5�S	���e��]��ݭ��(���\�}�gې���FQ[6�M|a8��[�)�oԑR�1ڵ7��g
����%s89��iM�3�ľ׹�
Yaⴿ�u_<�,�	q�_43��s��l��ب���'���1���(FNjYa�#���h�ncǤ�g��7D�^��-����;j�&�WQ�6�A�c�`����]Y�t�M��W�F(��ߍ6���'��.O(d�v��=#�'X�&��r��a'�����^)"|��**x��m�����-g�vH	o�ԑ`����i<H��7�!�.�J-�t�z�n�� �{���l�}Y��zD�~}|����Z�V���[K-ck/m������̼\�wh}�Ff����Rs�@���(.5c�A�t���/tֱ�D�g�JB� �+�KV	���v� ��F����rQg��O�ق�׾�:�6f$�u�W*�a��b>��y�4�am��#k!���Z��)��~�v�7�p*��Թ��j+�u��H��dQ�(᳃�g���$dI��X�;k�?n�S�l�]��'�l8�$JU�M���s|(�U�_���7B�ӝ�1��W�w�{�W�Y�!d�\5>�o371g}�I��9|>��z�W+|*�zo ����u�"@�ۧ�v�=O-�20�np̀�@D٠'M�q���~]W~�OB�ݣ�S�3�)����|6�Y�������K���T����L�
psF�[���4$&�`��%E��I~�W���ˣ4�|)�/1-E�r*��+?��$>qq�n߽�{���Z6�ǃ{'o4�S��dv�����B06V�s)�E(�����ۊ�YN^䃃+C$	�o�(x��`c%�������+Y��DeN�"0�/1lú��^z��c�
d@��P� %j�~��'1�Z���0�n-W�"�]G���`���z�F�ڰ��0��w�\�"w��tp�xf�Ln$$��Z��q���)7)��3RqR����%%��|.S-Q��z��*�[S�*5�	i�]�gx0;���ӳ
e�9#��%8�~}RQ�D�}���BB���@L!:�us�| /y#ias{�x�|���	WL�0�ISL���o9R��[.��_�sw��opD1倘�>B� ��sSi�vd�i���}�Ǔi�xc�W���f~xA9+]g��$��'�ZM���L��7�L��bvx,�F8��d#9�ܖK��<�7���تy-CØ�f���5M���`R5�&�@���'���:jδFG8U�ǒݺu�!Ȥ���49d�bA�yyP�-!���;�$�d���������5�h�GW� c>)�Q��3{n�v�jӹ��}�H�_nB
��G	$`��v3S��	���ȴ��VTT���s��˷$�QG�E�N��7�x.
��%&�j+((�	����~�ku[�q�߬���i��r�8�f��ӲjM�Ѝ��*Cl��ä5U�0�u\��[I&Ao8����伌���!�|惟м��I5h�!s��Ѳ�ݐ~�t�fNx\��ʭ}XL񱿀{N-�M���
�]�˙a��Z�R�F�sk��$�eúG�H��uM@�A�_~���g���!���Р�\��s��	�lU�;?;��8���dUD9ֳ~�,T��W�*M �$;w���h��S��f����֐�ط���]����#����1���ϟ�F�Y�a
8�`�����EE�#H��.bo�{��ޠ�[�����bl�/�|��1bm���ֆJ)��E"�-*��J6�u�Pq�1مiP���i�x�qE�۞�Sl��A��l����3 B�Q�.]�VK"�-���A�/�w�{Ӊ�y��j4O`��Qr�:�M�w��B3�C��w�{���u.A`�>��ί.�t����ٔh˦(3��>Ry�s��?Da2R�P2�����tDD��M|�]����;O���Vl�XM������8�ڶ�& �jT�g�&g,�z�k�ogm}�܌�Xl�ADs�"$��ǹ	>W~F,އ����Z{_i�|�oT-/����^ܥ<�7Fy���?$��#�֮O�ذN�sKT�/SC`�l��b��K9jf*D�f_����k�9�<jz�ϗ�P��rDs����"��F���Y�f?c���lϩ��`-���|£�nd���HR��V��G�0��C_������(���Ѐ��n��EQ�W�q���xO��'��$�"��/ >	,f��YO� !r����_�Z\�oos��	���u���2�9Z��`�W��w�Fy��K��F�e/u)Qd�����y��oh�/�A&��"�a.3{��~ے���K�:Y�C�-��R^(7[Hx{k�h�Q�Hcx��*0c�i�]�4���&��Ƭ[��B�g�[�C�_�����xˬSZ�Xa�'�f�RC�E~v'�'U��**Y�o�n�3���:�5���!!��������"Iz�o@!a���/u�̲���s�N4�4�1�k=�N���2�7�v�Dɠ6 \Hg�dD\�P��W�m	�}ǃy̢̦��8��珬�i��A���l�2Ժ��#D<����T�iϓQ-8�Vv{��it��{`��H�נ�7�N<���f��!7P�/�˰�!zY�vq7��X�Un�<UR2U4����f�7�j�r˩lL���Z^p>	�~�^>F��!z�`V4;����đ��Z8�"�[)����6`\|��h�|���)r�観V��,'+�^85.������������p����2+�l���+�G:-�Swؙ۸N����}�@�F@l���k�^��s"�rw���s~��rɴ�ݿ<�`��0��o���4)&��#W�K$�ݚ�����W; L!�]�&�4N.�[Tum�D^�D�PSG�zQ��d��D�;`�Z�]��6�~j���"���NI�X�����2p�_,����ܝ�<.��s���Ke��@�&w5LP��@���Npsf�٨9���"�;�%3=f]C�{ͫ3�5Nz�k�HԻˤ)����r�g$-!����rA���p9Z�{ )�X#b�Q�#_Z�x1s�P�EAZ�>d�J�TJ9"F$y猓��|1�L��BA�B����Y���s�=��d�K r�mL%�/Λͻ�|���tC
���xyyabcc#4.O��e*�Y��l# ;��<t��	o����v �
���"���Ŧ��� _���T�yQ䋆7�ݵ���\�m�ʳ�R`���!񿉬������p������^��Hjђ{�˭�l\�EqJ
-�vq9����j�>T�_m���%�2a��ER��i��]#ٸ��d[1Ѡ��Xt� �/1zn�X����OS[]�_�te�&�hMHk�}gӕ����ĺ��
���"}��_5�RT�����k}	���~�3�f+���.�Ҧ��=�?\�{X�ɲ�iQ���c�A�L_P��g����CQ�%n`/�fWC�F��J[�Y��m~L��9��R��A�j��u�so
ǚL���6U�'�y��#R��r�L� �G�E�LuEWit����̟W�x�j��p8:ڪd��yUnG�u�I���v��s؆�~zĭ5��.�+P
 �w�lK,����>��J�� �x�ʮ���/��n'��5抻!�
�M
L�p$�~��A�[j�O�d�E��j�Ѥ^NS�k3d;��p0�癵f����x]W�
[���;��,|`�\z;�f��Bs�J����_q6 �-�� $�a�&�_���y��s��	A)Y�Z���Bv�����1�5���y/E/+��ê������r�A[K�C|���{���Q*c=G�ԈWa0fL�8�K��G~�H4W?�$����^g�`F���V����{�g�cvG�և�fm��ֻ�&�b�M�X�k�#���
�ٮ>ܣﵕo1��57b��°)�@�|�B��n�#��`P7�F�c��u�9��Pe�ݯ��e��ۦ�3�l�1�z��le[����}��ڳk�Z��U���Bw��Q�#	 l�r��	-�p��� �22 ����aT�����"�c�՟uؘ�'�����խoJ�}/�m�%�8O�	x֯ʡdx+&�n�x�mL�7�*&��������I�C����=� �<�T���B(?}'p8��8��Aɋ:!�Lp�&���⫓乙n�WA [}y6�Rg�%�L�9d�8��Yݷ���\�e2��)9+S��TS�Φ7�ؙһh�
�qB��r���<��Q��巹g!K���{{��}�'p��)+N�&&C���)���*D'�%kn2F�������74H�8!b�.4�=В�h�]w3�Y_���56;��gE��'r���>1�UB�8�Ye���~rؽ��&�T�o��kcJa�J�a�s�>/cߓ�^����]~��-Jn�s�z-�è�L���/M���_f�Q��É�­�Uqav�Yt�.�o�!ߩ�g�R���N��~�X�W�B��h���ń:"��
�(�!�G�.n_�qhO��&~�ӏ*47��4D}0k�T#a�|aR�th���L6�hly1N��ŝ}I���x�՛}=O�R���}^��x��K�|�j{�$\>b�+�h̗�1���ǧ���@Ò�2�����v�����%����f�˅������U�c��`N�bo�k6P�'�	��p�XUwSJ�u�a]�O7w�q�M(�=F�9g9_��)!"v���V��Ӽ
Y.�G�%�B�N�᧓�U�m��<I��A!�љ�n:+;6��~x�PJʚ*��gR�������"�3	S%1�=�rh#��E�>��l�/����̋��M4k���;��C��9�Z�'�ᴬ�ޘ��v�L�E�����Єҍ����PˮX��7q���7̵7b��siBh���C�k	���`��70�}�Ee��s����k��l��6ON7V^�1��꣏P�s"|n��7X��v�p�+O��b�ɀwVp���~����c��N�Np�1Ϝ��I�Vjo�^7M�a�I���hވzB�!���\�������0���<A#�Dq�~�^��^U�s��\�3� 'd��ޕ�4(-�w�~DԴ�i`}��X�mh!�5֮g��t��B���'G���m�Ռ$oT���h�l�㸊y�*���8$7����*��"�.]�"�����"P/���7��4"]-j�>l=��6�^t��t��8j�U�\J;��\���%{��l�q&ki�s�\�v��펽�5�W���_|$N-*�n���S����-k��\�7�w
�J1�G�<|�-�)SU�W�)�5���2���!��i�+�}�p �j_�.pJpt�{��4�=	|8�f(���@�~��Gq�A�Z�K�l�O�VYMS�UXr���=�҄w�>��[ŉ�2?��5���k^���ѐ-|�A��s>n}��@4Q�*`ۢ�sP�w3�"Z���!�-{��)d��Frt7H�>��e��O3v�hk������5Ƕ<�z9���`��r�+{6W_�`���^�x~ϩ F�]��$�΋��|�<�r��Gw�����c���w
��Fx�X%aE���Z���1RƟ��9M	���p�(���@�etX�[�Tؓ_h�"7?{����|K��RL�Y��Y����'@�l�%q�`��V*�\c�bV��K��p�WO������&h�P�jD`V�ww����q�WOpF�L���*�[�=D�?�U��q;���d8�+�G��#f��ˮ��?�ٲ�&k��&�>�B����mY���۳c95k%�x�V�7]'RH{�J>�6��Q-Ҥ��ev�X�y�9�V9�.Ur��D�tx'�h��&��xY���'<-F{�zV���������'�	����B"5����(���hEˏI��&�p�䬑v�)\�\���o�p4�$oW�VX�o�N�����ˁ;��J�Yw�mQ�L>q��b�r����|��LOT�D�·WX�Y�w�P���t��9u�W�=�"0y/�@��jP;��G(��?V�@���̦~�k�5��"]$��������L��f��1;��>Յ�����-�_W�s�ABp����g34\��LG��׽���{�O���,:5�����#L���C�$�j��	�\��$���?�w@�B�N�z��g
$�R���E*����H@fp3_�[�^�KXGfv��l~oP�K��\xr�WK���'��%�v���˂7��Q�?�=�M��>� ��q�4
����;�pm��|/i��UqH��S�s"?��K�&A�85=�R���$�f�:��B�(��8��L��v�E��j������}�K�tbK	��g���،�`6��HP���Dv�iv;�"�x,@�V�g]���#�q�en��g3G��+Z0��4BI�H#�1Du?��Xz�]��관��W�������D�FO�L��rڙ���������P��H%�ح!��C�]����-S������ �����Meѡ���Za:�����J����{,���t�=�
�T�Ap��[,�3�����e�;��2�:�_��.N߾��8��������1ź��l����b���!l��e.�����#C~�!P�މ�u�!)����� ����a����	����7|���@�7�`��(dz�8~��Lݬ��l�z�BR�=���U�W?̃�@2�������*��qK�F�j�'J�]c-�\�O*!�c��g4iE:tS������u�K ,Z�,R��R��U��ֵ�lk���&< OY���_f���~&5�u���3�VEѸ�������8F���10���V�?׽��o��)�����<�,�c���?�~��7G�7�ͫ�����׭�h�^E%��x�t��k�H<؊�c�wX�9w׌jtd/�j��~��i�a}v�F5���)�P3�����,�-�����ғ{��:x	��� �t�SpG���°��y!� }�p>_TC�������r���؆�k���g7��XB����#\��u��%p��k�Q���F�"W���� տB�D;�h�޸�zU�fF��B�@-!�����'Ȇ�Ό1g��Ҟ`�S}���03�V�0��S�P�_#�t����3�S@���Q�0S���6��6�2�/�}|����/Tl�vD�"yӅ�����2"�Z�ٚ���.w[�ch��.��#<B�sjY����d��y{�_����8���d>^�<B%�ܴ�Vr�T��j����7*�1BS����4.޺��t�y��*���(�Y�� �(�h�`�V�86�Ti�B�zg����I�"h&�,��6�R�aNi�j�s6��ʙ6~u�Q5�x[-�U!�Q_pk�<Ox�j��T�qd���/�g^���I����ɚKXO&���#�"R��=��>�� []'��f#�W!���@���lްO}\ �qkB]�d!���+f�v�}���V&{�PZ��Mst�:u`�U�[�&w�/�[���;()��N5-�Q)r�3�F))�x�k������:g��"�nkC�2�v� ��y�U�����=�Y�Jޕ��ҙ�ܐ�rA���÷�Yq�����K╏`�f������\�#C�䔖����H��%mt��)����Xe:,�pd�h��h(��(��~� H�pv�]L�33�Y�Z����rAM��"[�/[d����#Inc�hā���|gp�`�)Lܶu�RtL)�ܩ���2���p<�d�a�.�2v�N���Y�3`��xn�ܸxN1c�C�p��?�	�u?Q|��r�4�X���M�Y����C�P��/"��t$T���O���tN]2p�0�Eȑ���3��f%�J��B�C<r�����J��zG��~���<���lN�� ��gĻ>��x�����8j��6�EO�%ON?�䤤�?��v�d�n-p$�����w�
�����V�h�p�q�W��m���5ڇ���腸�dY8��ؿSZ�_:`��A*)�������&f#�;\E�Y�z$�M/ժ�(Ed��W\|ԧt�Ԋ��M ���53<�������I�_�@��y
�[/&�V)%>�{�M�gs1zz�V���0�@Jzz.I"V׎'7k��g� _���Z�ȮE�/�}R�\��tn8Ʌ��t�F,�h�r��ǲ���iw�PWz>��=�� g``X�k�b>1�s]M�(_
#l@�T�� �(o��]Y<Y�4��3�_(�8+��@���Q���~�z�����-��4�/�(
@�1�}G������T鸆�Oڠ����)�nu�)��FLM����>(���r!����eP�>��b�up�4�@i̎����?i��WT��Z��b�y ����5�u�qJ;Y��72�8~����Y*;�ao������4��2��;(%yu��O<kz)rE�0KNx~�}~0%?�olV�d��?�lyF62Q^*��?���Q�;E�+JCEŐ�$�nwaٛy%�~m��:�3z� M����U�%����X��kM�e]�s~�_�$I���9bY����q�]��գ ��XeoY���巴�С͞���,��]1����c���!�ݱ����!
��`���N�����D��OfKΫ�����@�`�au\��X��=�	s��{	�"�3���r&���7�wDZ�x۵��.ՎX�9�%��vs�t�{#�{в���l�$C�p�JA���?����H��j_���~�]*���1�?��A0Ǐ��	���9  �A{/DD鱏�Ɖ�������2l�Ǎ���C��ճ�2��z�<F�.�B�F�O�3H#>�Ц�ZgV���5^�
*}Jx��F%D������q��m�������ui��ի ��A�G�V� 3
fL���Ke僑%��4���KD���N�}���ò/x��?]��2,��+�R�W-�C`k�]?Q�������R�\j����Qܦp%��y��OII�x=��w{����^ye��ŀ֦&QFH�3[%�Xp��lP(59��᷸���=g}�)&��g��ȩ̸��ݜ��*s��m���w�{��������f��]�2jE�����]AV����fSΏ�u�v�_s��{�ʶ�yp8����m(K]���l��ӝң�Űϟ��k뭇wNo���N�6��l�z��#�8�
�ه i���n@Z��^9�!�p�����K�-� nl"���7�HHw��`��Uw���� ��0��.��}p}Mι�7o���	:,$5��/�iY�v$��I$''k�9#0��*�/��Q.�P{�V����k!V�d�%��M�*uմ5�'1��x�DNi$����f>���}sR"��'6T�	gD38:��+t�Z��F�2s��0{��@�`�WV1.-�b����"�թ?hg������Yb�lY<q^r��
�ׯ_�z�֑¦jc޾=�u��M���*�⽋9�٥��C<�a���yS�c�҄m�(�g ��L�@��dRt��5r�q�u�^����^�q	(�(�]��{���(�F\��N&�T�e_$3�b�74�������-���cR��	U�z�ݦ�v,�o0�f>-�	�xR�^�M���\�t���[S{;��D���MXT9�p�iv�_T@Y���йa�bf��F.�}8�Ѝ�=ױ�;���T>M��g3�qj��&}���|�w'���_�	�)f�C�\�y&'�"&i���X�1/���i��3�-f���#����5�F��G��f5��(~mt+d$%}w$�+`f	硴�Z���V��%��1�(v�u��YP�K�y��lkr�*�*�d-�V��/�𰂴��j�97nYO����^!�'��kj}��QAN���E�F�E���1����!�wqi�V��je~2OYu)Hxo�}�¤��ŷ��������!�Re�֠�Z���3�r6a�_P���ؔ������gL��#�__n�hN�{���g�oi6�urA7>a.e+���`����3�g	Ŧ��-Nk���z]'������@(�7��s�:��&�ee5e7Ey�n�Ճ�cK�q�p�ׯ�\�Or�X"(W�H۬#��}�ssݎp�n����E9Y�h�N�����V���UA� I�����2�2R���'�e�E�&�d��FQ�p�����d�'�趹61��h����33��07aj�~E@s`S�.�	�P�6s�z'�D-Q'�;��+�$l�&(	��rC$撪K~��e�u�]�MQ��#A۵��+��m�/�Ƥb�H�y�M�] uyw�EZ�Z<<<�)zzz��P�0�#�F]bg<tC�p�̥t6������'׸=�Ln�La�!aq�z�g��C��w�A����rxԬ"� u��Q7H�7�[�i�|����4�D��p�?���}gdcC��QQ�9.���7� r�44V����,��>J�@��U
�s�{�R�����Ԓ[��uRۑV��T��A�H�-��D�lsXj��/��ߞ$��ꐳ��;�ɉ;/]�T���a͏�"�����A�a�����k��'~{�zO�����xqTp� �<ݺFޜ���X�Vl��g���aFz������������+qh��?YtJ�	9-�3�-n2���"ܵ��uP�jֱ�+�zEc���pVn�g�trM�}��GLL�e?�;2C�����B?`�#w/6]�w!�Cԥ,M�/�������թ^�W�����K���n)��]�Y��M5��/lY�������d�~���Ƒ �2�'�X��/|X!:y��]o�j�B��к�}'�M�oN�7���ЭE���ԟ�@��[�/��Dpb��\Srp(4j�����*�&d?�ş�^x9##��K 2I))���E:').S��G�XE�,=�7�(תU����~h��$�����G\���-"�ަ18G)���I���~d��U�è���KR+�؀ě=����y��O��I6�Hwz���/�#�{"�bzVN�N��U/NQ��/��-�g��	�_�U,y��W�d\��o����{{�M�x�[A�7B�s^�h�3�7C��Z�dC�Y�gF�N��'�Y&�4�ןX\X�����_����W���lr���\�vdz8Y�jP�f��O�kSf�;�	����:q���Q��I�QU���UEC#�v@QQ���AZhI��xjY�`O&�2��?{��p;m��y�CM#�����|��4e2�����^�31��2<�8On��1�D������K>���LX�?ҀqAf�_�a�\		�1l��e�@Q1ز�Б�J�t3tky�g����dB���"���lb��Jl��}�/��]��1pO�i�ה�f�n5I���E}@����������=B��'`@b! ���Qv��qXx��������2�Ϋ/'L�}	(
^Ԟ�nt�/�|a�<����566��N	TRR2W��=M9U����k��������P�ۥ[���I(�\��3�ld�%�u���D�!��_]�[�Z����ʌ�^����R��{�.�{��.�|���{1�Ἦŏ#?~�	�M��r�ʮ�{M6`hyu��ܭ�~���,Z�ǰ��

h��p��A������۞kS��������ZJ�pDf�!PL�!����5��1��Z��ߔEf�fv�'n�>�wo���}�M,-<��
0�>���n|�;܏��������"� H;r5%��ψ��%��f�����C��*V��23e�ׯ�JKKo,�k���ʹD&RX�;� ��bq��M�b�`��5�f�����f3�f�_f�m��׎z_�>�*2��h�NPK�u�q;"�7�os[g�)Ʃ���7����|P\�/+�bcc��=��}�Q���	��\G��4����C��p��!2��i�bgE�[W}(R�����\�C�YF�*@Z��^����w���[�xV��R	9���-=�Q���Z.]d���h��}Qp:��赏��t5!;�7mL-\�"ؓ�<�eg�����7�?��ؓ.o��ƥ�\ (�=�q����{�x��Y|ϫp��L��|	]o��b^�����8�)��3��uM,�Y��$��_.M�x�&Ĳ$.����񾧙o�4��~Tl3��kW=u=ww�z�o�E_DH_#�7y���Dٺ�V�*��Z���k�
��Iq:  ��&ʷG��h��QH�e��1�G޼��<��:QP�HE���*�����ӱA��蟱�G�g%
�'W�i�PP`�[�K��zkwC�����U} YzV��R.��t�O�ƍ�!i��R�� �B3t����3b��m?T�mױ���^;Z]Ī�5�a���)H�u��rw�Jr{�7��m/gQX�u"��Fdi�7�\>=b�����]l�QV?E:�Ѧg����Yh��xlL��p>�
��3E.zc>5^0\���:��ɰiZwJ�k���˻lN�Ї~O����JMI���r}X�`Jж�9�
��� 9O�ܓ�sޫ'�^}�������w��'�1���/j�:,�4��%
�;�ߝ�������3�Q�|��Ȥf���fU"����e�8�V8,S��<f}�***pR��!K�� �(���r8y�NT}�4O���yW��-&��i~r?+�E�%���tn�6�sg@��Wf�U�@��ɕpX&[��fF��+�Gg��gZMH�:y} �y� ���'��&�%���۔q�
�۩��A4�Uj��^�a��̽{�O� ��\P��M��P4�"g�垿����v��f�����/�������epo�vJ�0@�:���hw��O�x��nl���J���q�)�+TX����v+p^H"��~�{�M���8P �}�Ƞ��� ��22 m�K���7WP�;��~q�OT�F����.�幘���*�0�h;J��f�&?ۜ7�v�=�T�7jU�щ���K��K�0uп#Vf�{��nA:�� �|�xǃ����Oag����!V�������T55�w�g���RhF�k	���W*zH00�6��3���m�Cn}M��j�_҆D4��p�X-
DDM���Gr��~� 0K�����f��P`�B/�;��s T������Oϊ����s�5X4�z#�����P���{�]7��r~��"d�!/���v��'UT�r��а��� tT�O�t�|S�AB2���P����<��`�Ll��;���3�u�>f^ĳN��<$š�]���Vp>bU��:����3��W�c[��׾
+���b�zr㯊�8S��^[���c�q^?�^�D�|'��r4^�F�ٳ$�y�������y�v1�<"֦-�[s|!>nʆ�F���V�ٸ��%���v$� ��Jwϛ��[��Z�:8����[��dh`��	I|�O�����8��c��C�%�kB&��H���d�7Hn�Ə�.�T��cK�Yw"5P���*��iQ|���.��D�!����i���2�ں����QA�Ư*��T�#m՗�o������C���kG̠����k�°�So	n��/Թ3e��9=6���� גד���RA
uΈ%	��}Z[_�jnoi�)D�.���#��
�$��hs���:�mѐ���,(@!w�&�'ܼ?�A��Q��.ߨs�����W1�u�Ɇ�SY�/�)�����4�b���"?	vk�Z%Ha�Ι*�_�(����:��B;@$rONi��Lzr9�j�<�������U,8eF$"ep>�﹟��^AD%c�1P����QS��И�̹9���7�"��8���Ȝņ�Cu�����!px���h�O�����刱���bk�>9$��̥��	�!����sW�h�}I���W����E�T6du�,Vf��Q��aH�vx܂0���ԝz�fo1���dš4WF�� ���p�*�ۖ�MN��],i.�K��|�ռ��ĝ9gPN��s���k�Ͻ$����q��|���i��-J�zڏڠ ���2�AQ+O-�"��\����~� ���~��*���!Qͦ�i���*�_�)tЋ��m��1J'%]�s �p7�Q�zϽl����g���	����X��E�7}hV\m�C�l��㬿��۠'-Imߤ�Ct�n�|�\Á|�_��v�o��_yXhe��W��g�U�Ф���;��e�J�����!r4�t��ƧN0߹� q/�3����᫺��i��V)�t[RZ�Q�j̓O���椽�{��T�]u�U��%���~����pl�cU��ϙK��%�9��4�*˕V;�ⓀE=�Fq�}��>���p���B�~��2n�$V���G�ڰd�'��)Q��1t���� ��uC��٨��X�8~�wY�Mewz��S�����",GψXlg�ϑ�E�m �IOaBh��6��|Q�)LY����]|��&~��C\�<�D7i�M���^�$��@7�e����z;��/����O��FC��ȴ�+2��F����_��ԯ�z�Mp.���w\�2�Y|��jzD�����N��n�b���Z�u��N${/uSm�gP��v����t
�1F�V+���8����)���;�b�S?[��ɡC���;��.~���Z��b$ۅ����|U�����t����Yk3[_�˗n�j�~/Ց&�0]m�ﰈ0���{vş�������j\u^����w�����E�l�TOr�����j WQ�J��0`fS�������/_��R������,��p�_N���|��b��kh�������C������6����i���G�
d͗�����%�]Rr>aUu�^$ ����H��[���Qv�{{��~���������t�d�g��Pq�����{5���^��� ��NS����k�%����qX
����C�Ti��E�㥝o��y�%;77�0���r[TC��n��20����2/UW�M�8*��y��sl�') 
<N�ω�n�Ba��$]�,��Źү�hVW}(�z4� ��7,}'I�\$���D�Ztz�>�k�A�,���=\�dn�ݤh��0ᐻ�!|~�؁��v��"����8�׭c����R�Y|��;R��̥�f�_!�o��#�;l^m!�q�V�c=C�d�i�S��2:H/`{����G�cs�~fn��l�c���y�?����d�u���Uz�u�۫0�e�
�R�k='*�M��&jt�(R�f�0�g��=�^~��)i����=	l&�%�H��;�f5V!-'������X������/,,�3����ohH#�3��v���{��%w�I�(��j��P�qf w�/����K�.�]�]�v��!�x����!������LV�8�gbf+�I�����;>+��	� �%�jTUT�0'�|/�0K��A��S��C�AE������Jir��%�����ɦ[9��sҾu����j�7ll�K_��^�]y#B�m�z�	o���S���]���z\��7��cQ��[�N�c�^�����rӪ��XX
O�g�P)<H�b옰�e�ͽ��������>�k7�������P��e(_{��Ǖ7,�{.`�������y؉��$G�y/L��U�k�?�>C�&�%�]�¸s�Ŷ�=�U4�r�"且{*��OS�r�K��j�<�2aH�¦V����[�X�
7z��\}�+�`�&(�t�<�řJ��N�/��������Yq�.8�nu[��߲+j+�I����X�ogd�P�_�6`?�}�{ ������K���`���y,DJ֜oq��{�l����OyNֽ�HQ�B�;]�0x�ďm���(��d_���[��E�q�x��A ��p���V��4<m ]x���X^�*��:BIr#��m̄�J�Q0L5�p�z8�^ک>�=(0�Ɩ�F?q&k�f�{�,ܔ����=���iXb�[<j��*�T
U��E:�K�G�zw^��M�wv�]�g�?��{ltJ
ڿ'��+�w��`Ju�ы!�(Ps�"A�c۪q�ϕ#Ï}(R��!�.�w OX�x|���X�������H��g*Z�M�|k��fH�ڳ�`J���]���>wK��h�v���BfaȯN�����V{�_�x�ܒ:�r)�)����c����\T]ٲf�]0Y�s�{��w߇�B̵�֩��P�!9Å}�ұ�3���(�/���2^	��Cٝ�:(G@ϾR
�?�*[�=m�ܖ��Z�����Ĝ��F�jTwxJAh�>{sQ�o�y�}ZW{�����7$dqi+})�JS)ȒUPڣ�
��m�ǉ�+(�0�(n}�|o|�]f�h�f{�ۨc�͉L���񺨠KW�I[pCcT��[&~�#�pz�G��8��a�n�[ ɐ�����?!Bn�X�\�߳G5-�a��4�jB�j���;����c���Ⱦv pW���
v�8�qSs����[�}Y���Ƨ}��R2��:	��S47���	��]��SW�ϟ#���T6��{�@
;�C/�:F�RA��Lm�K}M{�<yɐ�_'<�`ʡ��T�����|�$�^UӟB$*��(�a�����Wa4��B��⛛	�N��2�V�Uȍ�1郌@;|�i����]����������\���C�d
L�ޔm�q���e'fs����@����71�=�^�"Ç	>���v��ea��<�j��=�yl�a{|(���:RA۩������mB+؁��6-΋4� ��8z�@�Mzi����O�|��$l�π�nm�&���#ãs���X5	��g���F�Hdpm������QQ-M����P�
T$�H0$�!�J�!0dQI2� 99�EAD@�(��(0���F��������<kݬ�:�C�����UW���]g=�1i�^������ᤕk��&f�잭֦f:�lL���[j�	�4%���2'&gʖ̫�+�))�uQm4�u�Z��-��i�9�A)F؉@�k�l#0 �YH��?ұ�YE�n�b�� �y.~��q�/���~Cg�j�[�3z�5���]�,�g	/��Y�����ߔ�<���7ا־����/(�k<k��y���R:�]P����p�Ƥv܋��:ܘ�)3�j����bv�-�tL�'y���27�ޅ��٣eKzP�+��;���#�Q3��0��g[��TqoPz��L�l�L4(˱q'�kL"��C\ۖ�b�7U�Na�n[Xv�&�J�A\h]�^���ゔ?�\���:<�b����Y������B��o�;�r=]�tl?v8����$������}�Э�S�?�%��_i R&�i,frʨ��p����h�.�F^>A��1���"�i�P�o�)���Єm��[F����q��s���O]-I�^3�Y�{<sU��C(e��?�'��������?��5ieV$[�J�N�ޯ	8��;���@P������y���]B�PdS��A�Or�+b��g� ���Ͼi�vMR��K�ƌA���g���^O�
��Ϙ�<��s��Hf���I��;���Jd
�$��A9��w?9|Fk��,��n���Tsd<�p��c��q[#"(F�B9�n~�H���#2�i����%-e�>G�<6�N��iI��&�	��b~�/	�)f�������Y3��֯�(�M�5�
��+����}������{���uOJ-������|s<�ʆ!RAe�vj�Y�#�S�o^ϖ.w�����W�5i��^��}Yk��n[�݌|����4�6x۷w�:�/mԤ��/�#��[�2�w2��q8�%�&p�Q쮢�_�en.�2����	�%�p! X�<+̣����d���薏�t��sػs��/z�C1�>P=���o�h��2�"W`��0c�
:�
"�N�1����~m�3�f��K\�:�`̓�Z���3��3��P:䏤@��q������U`X:�� �?|$���s3Z�Ν��MR�DZ:�ŋ��-�@21)����vss��Q}��ܾ�T^^^MK+EIb�V}�U#��)�m�M�P�GAd ����$�GȕZ��L���>_y��!>?�~&[[{ۙ�)]�����$m�SOM�Jĕ=��&1kio�[�v��Ko�z��@fӓ@�Ͻ�Q��Zb��P��W�$��m�}����`�Q��2Q8��X�$Z�����k,x����|m���k��"����qu�Mf��]Yh״�c>����y����������~_%�v�����Ͳ4�t�+Oxs|)kb���F�a»�Ɋ�0	[/C-q4�[�$xݫ58,�V>X�$>C���p���ii���<�Ozc7�0�_A��ƱmO� `�����r�0��b(��f�A���=����'����_bxj�U�3�Dј��4��\e<�_P��u* �ajv�n���*��x�d�9߂n��Hl�����h�������C�89[D�0QM#5\�C�����&�%:)�`~��_��wCœ��)��fl��]/��;�OCs{�ͽY�f���ʮ���o��8�
[�o�#яq�%��6���d)��n�}�t�Ԥ��()W!r�Dt��7]����e�sGx�흾=�G���Fַ��������g�3�X���'2 {��Iĝ/˕9��96Ȩ��p�!KG�G�âd6 ��w2n���`'7Z���b{;}ewM�'��e�d� �J�eM���,��b�������s�_ƹ�(� D��q\5���&{z�Ao��%OI-KO|;�t�:PVE��S,�p8���	�	�?.΂������g�hB
#�}�(v�-q$m�%Cƞﴽ}S�&�;�S��W���/ �P�h�+�+q��an�
o���#7_��q���I��F�͘ƭ��4x��.����E��&�X�J��)�,Қ
]���ef�/ -�Y|hz�g
��2��JrW�;~&�V�D���QN��#��6�?����]z�i�ι��<ĉ4	귴_b���~��������d�k|�n�&�_�N:�|�Q�IC˶���ŀ@�{�ǖģ�g�т��};�A����'�%�7���S����9��[���R [�d1�~����vf���n�� ��^�9�p�@�"���nr����c?�Կ�c�����@��fB���-�s��׉���x�t�6�Q�d��q���j�J�b���5
{^��KQ��̾��	�
���ͿC=fR�?�'j�O�e�K"J��:;��o����]����`'0��ZBZ>FCR4$���w�7\��V�{uN"�����"}z�&���<��edG-�ɾC*-�9�)�-c&��E��>6�fHh��8�еfK. YD�Y���Pb����-�˲�{e��v6y%�E�Ѣ�O�D2d3]�fVZ��x!�Nw,�؊W81�#��[� FbX�*��M-������V�S�����[���0���N�j>"m	���YS�����ٿJ�rY@^3 }�A}[ҥ�E4<56L�X��
�:��_=¢}؂n����WP�FG�Ji��F��,?c��lI/�2
V �:��U!M@mI�S_<Ew�,n5S8���v
�E���(��tY٤[����OS����v�Q*t�F��qh让�f����T������2Qi�4�ט~O�M����MR~�b��4wՔԽkD�g�{�����ӓ���t���:��]D�k���BQ��c6k��A0��h������U4����X֤��{�n�Ά��>����U[�y�����)�@�ZG㠋�,}����@u���߫���Y�%ɝR��Db��Z��7fȁ�(L�"d���8 ��@�]�@9=���&i��$�������;�v���~|p��Hq�
]��?u3��eT)o���L��k�Ή���E���k��Uݱ���5�AZm7}��Lj_׈�N��?)�Ä-6$wr��f�Oh��Trѫ��[��F�:
\�|��*�;�Q�1W?-�h��u4 5����2V�	�PìV�A����}}�� }���I9D^��2-�}�\a]�T(�\���c�$\��skuU���ꃎ��F�J�V����2|�A��vi"�6��/�����$}ئ�C\�H�!���1tII��b3��j"�]q~"����,��,�^c}�2���� �}t2�WV�NXm�î2)6���p�3aV7�-Eģ��_V�*~�j�m� �㏱�[�Nc�P���dğ���0���U<�[q������	�t��7��A��C�t�jL|pp�l�1�H���nd���n�~���~��#-�d��t�XPӗ�G����l�	��q�"��J�J�&pD��؆�ff=�G�iQ{Ơe�i���_�P �,�S�	����Β�,=4Um����	�S�r�;Ǟz'��W��)l!����޺
t���D��*p%�CAu�⥿��,�����oJ��x����b���:�E����`���W�%u�}�DO���ֵ9
�>�Yioމ^v�{�>����=B����v���KQ�?E(����u�n�h��υ��Я��h�B���5��Ao�w:��[~�"�. so���OS�퇻�89�O�5\޳�ڷFa��g��GO�����n����dtZ-����e�����R��������bH��G�Mu�Z׫��S��)�Y2;�k��������]�qDt4����i�(f��f���N�[k��b��d��M��	�7A�eEW��m�����w����o��v���D���H��#���٪�o������p[r4pr���=��mjkn���R^��>�7׵��mܿ킽�|�O�VJ��w�����]B� ��o�o�+mN��◒����5L�Z��23�r��Y&Ž�wMI.7��fe�%$ZFNWh���5�`S�X��UgGR�p�.�>�&kzU���s:v5�A�0=��0�'��ym��s4��jsnk��C[�����K�U�/����c�i����)N�$��깟)Z�0Q(��<W����S�9w�l�9�{	4_��:3����ۘ�5��Pة{�ў5�b�䧟�}j��d}�{>���>��I\BR�7�U$�b<VW8Z��[yյk�ȥn���s
�j�QI���O�G��iC
WQ����8�0u���9o3y�l�b��fz�W��)��WǬ��<Xyjr&�xrV�e��WN����Z��������$F2�O�x��پ��Ԕ')�*C���U��v�M�dͪy.,��|�&��c�Cx�Ȣ9ٞ'��{�:��Ȫ+YS�β���x
ukI���k�2�r�MS�c{�����`��y�iO���X	�9�'%dyn�r����r~��۷�3���Hీ�tjjq	$L�l����.���l��܋(�{�:lL?ʲ�ܞEn���I2*���UX���E]�S�$�s��p�ۣ�{z�929H�+�r���W]f�_�*�9=\Ǧ¯��D`��W8��9�<4��"D�y���(L�l>�{aI�_�8��_��7j�)4�H��)�0�t��Th�V�#��{X79�EӨi��(|����Q8賥�7<[�!��B����9�]�"dK�$��<1@79X���j�q��u��f�{`Nm1%�!�JVL��c���*��Y�K��b'g�6I�v�Jx�)uEV���ӆ����^���T�D����"�8��U����<P�<9���U�(x��*FEuCfvNA'1w�����x�ٞ�<��Y��jIct���g�.)p�ߎ�R�;��g�F�����"�<f��:x��N~�V�p۰%w����!$��> �Y�-�r��2Y3"ϓ��lg[HM`�S�f��>��"rY t��W�=���)'������������O����J6:�j6��A�b��sf�	Յ������p}�̤����}z�V#z��5��}�<�
r~���fE	��H��l}f����}C����q�e�W�OJ(�����(�Z�����(�3�r��l�}9v�����T�{����q�UTL%��lR摂�9���Gy9j��zĞ�ON,"/���<�z=E.�����e�L�Mu��/<�Ű����(��j�8�ŷ�*�y��C˴���50J�E$��U��+�q	�y\���^�/v��iz1P����5��(��|;�E*\��I��0�En�������E����:���+rQߌjM0'���X��sپ>w'������PUIf��ꗕ�Y�W�^&9�>̠�̭N~X�W�'k!���»�l���0Mv{�xP�5���J��<�&��:;/W�|ɍ��=��r-f �z@˕�����/n呛����ց�@�G��>��W}�d8ᶗ�b�h��H!�r���T�H_��.~r��Lyb��y񂱁��s���}hɞ��Ly��ѹWc���U������j��V�����1���)� �C�{�P�Q�59]�����rO�b@��@N`��&9�	�J�d[*8���U*��#���h9 �I�8���B�=}ӈ�������]8�r�[�(;���V���������x.ߕ�&���
ƃ���S��;�ÇA�o��{¾�7�yp�[Q��r	������ޥ��lNNXu ����fmP�V�^����e�@���%'������6�����W�/-!�2�NW��ߌw�8'O�`��:�z�N�z�F�AE����13���"	x�ĔY� e���ɮ���+Ǐ��>T��/k��u��	��..._��[�����3��:��nȮ.8���=�����Ns O�ued��	r��?�nǨ&�I{�v�AH/�� m��@�R�'�[��]�1s]D
2�bd�p�6�Ǌ��5d|��\.��ߐ�����>��CE��uJ=?�No���h��n�IkV]���O\h���v����t�2�J�1;,�:�sss���"�Z��BC��L�;�R���D����8��8/q�_�f+VR4��-��hNer���fG�~���tbCתc���?�6�Ѭ�(Y�a.������ �I���ZY��ہk����u˴5���qgn>��z�Q\srB���'5˰��x��m��6�)J�y}��W1
��ڌ�{.�,����Ö7֓�)���1�v,��&
L�p����y`�B���U|�p��)��\�s�oU�\%���შ��r��ϋ��F]��"9�',����$8�=q"	�����y�����K�"������h2u
��5��1�6�y,��\<]:����sc����;v�d0�v�x�n�!$�
HR��A_*o�Y�7��ɻQP��Jb�Pb6Mk|�`y�Sm+�|r���۬bوZ!7�l�|�~���jk�Z�4-!�0�N�ufV��<i���1V=A�	��2�3���C��@�y���\4Q��q��Q�i�DP��)q���)l��"+��:�����:��ʫ�웱\
�)V���4W,������U==���0������U����U�Ӕ��O���0A}���?[6����b���}�t��Qc\��D�]^M���憕�����#��߻��d���Rɟyã#���Rȶ,a
�_Ͳ����T�;�P�)�4~�l�E�� 껓��!.�tg�24)�y?X�K�����^��ˢ����0�C>�?u���[��0���:�͙��$�<�;o���d\3��:S������ï�z��/�W�9�-��@��ɑ׀���u� T��6uD��
�u�F;e��	e���7u@=<**��;�288�ʡױ�KNo��	7��z �lY	��d�Q�5�0��r����4�^(v�f�[>������>�Fاϟ�3��T�N���=�Ɔ]�sU�X%�!�����hX:���bJW�X7Nk�\��K��ޮ��+�
L�Rz=%��p���N {�[\�)���Ѷ|3U���<HH��6	8�n {7����^���QG����g]�0�	y��[	tڒj�Ee�0k�܍��.��|�9!��{�n�����4�k-{��Q��3�@) �5zr��#�g���s�l��(�7s��b�}}���}O���g�|7$;��f��f���Zv��0�;Ǳ�����ܾ}['�K�q�H��ϳ?uQXB
��Ȱ��C��ȳ�.��9�p�h���Ӑ�fJ>�O��C���e&�.�t�l�\��J�u�e�9��� � �k0�a�q�%�r��T侀R��m�ENe�-�_���������2s�t"Dt��p�c��Oc~���S��-5��YE�RJ�~=ٹ�2�3X���f�	�Jg|t,�U��x[�T^��@��� )v�MV�:� 6ճ�r !Q6
��4�Z��� ���Lo�6��x�	V��}u!q�A���zu<�q��4RY[����(��� ���2m�)-�&�Te��U�w̎��t�s���V�=ُ��x�ha!�0t�]���PF�=�%5M���e.�Iؘ��nu�T� �O���N�&&��UG�}�,��h�q4����>���,�*���:u�Tᄚ\S���&�)!���z�F� X��~<X "�_�#Sfωw�+O�<~�W-�vJ/� v��o(��a
{�no�c�P#�;s��s�u�������
�0(��>T�`�z�U��3Uk�+;O��e�#� ~���`I������m�{��XyD�T� ��ӗvC�"�Xcݗ/�ӳ���ʵ4�
�{�q��i��|���z���;Z� �SBC2拤<|��|����X�#�D��U�T�
��X�Y�R8�0��E���A"�䝯�`b�!����������G;�{#U՜C�k�M_�Fg���pԡ�����p	(Z�܃�a��� �%>L2�('�������I!��o�#�����S]y2O�>�Σ��O���)�w >�����ɭ�y|���������,#��T��~���c O =f3}e�����ڐ3�ui�d2�>�Ģ�S��!$�7���{m1�rh�{�i�"�EK�3�"A$Uei�̌�/ޕ��]���^N��&l_sH�g9d4�F�:� ?����E#�v��Y[�P�?g��u�����D��9�t�#|*7>s	�[�p:A'b��؀��ƒ��T��]�~t+�(��OE/��\�r�5��|���e?!��ɮ<�/�����mp3��~��sq�A�5B������=g%�����P�*`v�A\�,����z-p��+\��]�6�m���_ �}�>�k��3�&Ú`�9-����q��YyG���-������~��JQ�OS�7�I/~��J��
[��@��"A��0~�/͵��Pko�L!�"�ۄS�"��u�08=��o	��@�A�Ev�GYȕ�
�b4g�AJeJ��=�rҵQN~*�6cx�h��k�sN�7�ߟe���]+Zwy�#�M\�Ph%^������?W%�C�B
-`�s'd5�~��b��}0���q��Z8���� �cߠAv0��B<��e�\!�*<=�]�111Y"�n�Z���h�Y+���Hc��R����?�F8��3~����z�=pi���f�7 b�Ed�?T�)��a(T�%��6Lpz3�Y�����d���{-)B-R���� #S���@��}şC8d~���u�y==z��Ri���L�
;$w�>�y�:�5%�}z��ץ�s�V̻R��/�N�\�x���im���"���������_]&1��1n-Z�o3*��s�
a��K�.a��}�j�Ϡϟ?����]�l�����4u��jrO����Aln8��<f���<��=���n��*�$��Ⴌ�J�* å�kN��T��&1�O��	{�Ί����u������ B(������sR��E������fSY�u�t�.�w����3�;��n������U�aPyN؏���E����s�*/�_�}tE����+n%�t�̀�����i!Q7}�NՑ�< �	��V�dmF߿��.���֝ս%/���d��!�-�F���?5m�?U��U�ͽ�츬
������D!�qV��##oM��)�K�.Ule2	}ۈ�f��/�m�8�~¬��'��J[t`��g�P��k7-�����^�)A���s����_r5���	 ������|5t[38�s�P��n8=�t)��A���˗�y���З-�(��[���]��o,��}�P�;e-���I�ى�s�
�G�LE׻��9���&�QI�z�'m�G�9�{��k�_�x��U�3�c�U�bgu�`?4��aO�_��Pc��[ӕpu��$0� G�b��)�;S��x���Kf���xӗ�P�[��7aK�

�/���V�?|�w��Ab}����N�D�ԟc����o�b�׹�8ޒ�""����l�����:0z�8rq�4/o8�HJ�#���G3��Vr6�����>�ϝ{ׯ{st�wh���-�(��QP�	���~t��n�W�g�\Gxx8��h�`gMoz�Uy�W�
�~������v�+�3N�Yo�$�h�OP�j�RB�ë>XR�_DJd��<~)��24�Gy��F��'��;�m�}�x����D�H׸ ]����S�{�R6Xr�X� �d�>c&��`T�q/*VF�B�pPz:x3`p������=.��6����X?;v��M�����7Lq��Aߏ�9��O�xA�0N��^���:3�2��]0�_�J���1/_�ʽ��n�`���J'������p�}��˂�������z���	5�DS�/o�R�P�a�S_G'͗�C��v�ί6�/�/��K'�`b¿̘(S9A~�DhbDk��5��TA�4`����� �T\�h^M}N@ۂ<���% `� �˷��R�\~22�4:�b>z�fP��t��,��l�� ��d�˷fm:pk��ܹ�U> ?�� �����#')�˫`\��d�Q5�#��ӿ�3焄Գ�#KPS�M�v�l���/JM���/^�Xq4�пk.���n�+�I��3<��m3�������v 9�j��8k�y����iW���VG�Z�0����<	��<p���s�U�(�^^����I`������A!��@���	��i�L�i�Y�9��""�S6��q0T��rw�y񙺚����ӽ��q��wpM�4k�DJ
�������$���!RHDH�ف���6�@�a1M�W"�iP����V��cgϪ	dNOH�EM���	񁏭�T�Z���4W]�'�ɺ�/�-o�Ű��,j�$ps��K,"�X���������w���R^���e���Qr�m�����.N5	�C�j*���%c���yII��������|T#K?��I�� 
�/ٲ��"���8Q�j�z\���V�+z��R���=�or��<w8ؘ�r�
E�R�X���؈� K"R½ ��,�QH��
�E҈�`Uɤrt������?���,jk�e�0lzD �/>$:�k��GE�:�y�y��]ePر�c��U�O���}������t�}0�A���`��[\�ub�Q�ۜP��֦�D�`�/|W��ס,M��' ��� �&���ks`֕"���K�Y��?����$V$�&k��r�r����U���	��}>���� '��y�{E/Vz���`)��2��e�r?��2on8�s� F]O'�=�,��chh�X�[�,�R���>��:�S�^iW��;̘�����+nLmF����C�	Pa"5�������%��4ɲWd��k��ud�����DZ������"�}kS>.+��j�m��9sr���6f���A��<�kA���g��@�i����L��`����N^��&�ݿK#�i�2��D+~�e[�B攔�/vF�O5r��/�TNh��V��$o�4.���|g##<�`A�mA�zizjݽ�Z��Y&2Ik�@-�y/�@���?�s�>��E2-��w���&�;L�gY~O���^d�Ee��k�$�
�K]������Z�2�e��2ʥ�*��@\�k�� �D�AW�(*
��`�JJ�� AGQ`k��tž.�Kz�U�Ѐ�kdV���1��f�Ў(X��� �_)���E��BC�TPQ��+ =�E}'s:�߄��$RL�ڍdm4�V��x�q1r�s3�T���ʆ�����T�h�k�.:���.?ᨣ�|Cۤ����de��M(JT���P�����לj��zQC�o+~z��k=��=dIC��M��ҹ�+��)�h�Gv��u�OI�K�>�\����`z�dZ���NW�Ȣ�;5��ƅj��~�:�Ț����p}��p
�Q��2�dY+�3����:����K��s72��Y�t�&�f��ļ�*�D*(�-�ԑ"-�Wą�S9�ԇ�n~�֫Ӈ���Q���<�[���8	���������0������� �+Y������.���+i]��W**Q����������x�������J>���m�E�R��O$�n^'�:��L���' ��1��]&"����h��'��L6��?{�m)��Т��Om��[�d�yM����?�6��Fji��ܹE���hbj2K}����R��n��}U��� ��|�0�(������+~:n����V�eM�)�
��)&�t��6�*X�=*����W�[���T(�i�C�u��O8�����]U�Z��P����,�3��fc���KV�?�aUԛ�֦&3���A��fO�l�2���j/�`���6����#(�!!u?���_��?����A�휄����b�3�t8d�D1� ��/���w�U�nY@��8HQ�(��,1Ns��!nU.���؇�p�Ic�ص� 	b�j�`��@���X5ۥ��|�� ]}g7l�������ȑ"�%����A�7t���;7B5���G4|�MUi<-k���7.Q�"�e��b��M*"��X�ȟf�X�J���Z�	~6�;�%����;�}5����Ú����������2�Z`�߷�rޓª�>V��4h%�M�@�g��|�Պc^kA������%�P,g0�܍:^��&�}BZ[�q��/CC���3�w1����,'#�=��6��y�O1���N��Z�?�����>�c�p/~�И��Gs@rc�7-*��l�:j���.���W�/2%�VO�3o�:�~�4�8/!'�0�M 2��=�����먝#L�?���O��b֋� '|g�Z����)�gc���q���y�z..�:o٠c×�=�H,kܥfn����"���x3R�TqP�b���� �6�L)e�h�'D����UС�Zd��R�r��d������Ĥ>�G�M�|�����+���#�	�8�2�PY�|y��p?�%�� ����.c�c�0[�)��p��G�5nJx�r}l�J{�;��vQ ��J����1��Xu[V�"�^�B�?p�2������@.����*-���^3��.kU�Ըn�=%&����ז�q7�"F����}+U�X]���Vjtc���4�44��\K��:%��9=u�S D4\���s������Gc6��@��etmz��P���3�Ū�a�1.�M���-���� �X�zߕ��#����CM���{�X���k{�$�j������e�Ef�bG�}����om�tC##�����5���P�L�X��g��&��[R2�4(�A~H�x{����S�,�~�9j
'�j��^"�:O�pv(3i⡻�������v�[�W[���,!�j���յ�ik�+��= ^��DǭJ������+A?�W�Nsqq���A��Ϋ&�v`��-t/^`�qy
�;��VXӘ:@(<�X̧J��99d��<_���3e��󤃇�rf�Bf��A�]\��"��~�|���Ħ�=� ��sM~���!I�us|)q"zz�ܷڢ�����L���!���7&�T�V�u�NO}}'���NJ~��ɼ~~9��ˉŷ�#��\��]Λ��ݘ_u�(�`�6g�KO��}���Z��c{'編i�&I=ECAk9̍��ݻl:Ϸ����hK��1�i C7�ނ�BtG �r=������d���L�īr<
�g{ކOb]1�~fEj�~���& �qb/���A�J����/��o黯-�A�
��|(�e�]�h,�t�����7��T�Ůj }6ny�����r:���9�=p�w���Tco��F�mOpC���Ĵ~rM�d ����iM�G��,�<�Ƈ�w�Qb�A�S�7��Cxn�"%=�?V7�k�w]��z����$=;�O��X�����?����S��GܩHcJ��cpS�%ī����gf�-���үȜ)�ԕ���(�d�����1��j�t�+f=޵�d!ݣ=������͔L���'2��9D1]��tWI�c'�
�¶��ʰ�`mE�b�\��)�"�����+P�!�#Т!Ei3���
͈a�����jY�M�����0�*m��Its��<K=PH��B�v��e�x�ngG�u�LgIE�!*���lxkC�(���9CQЧ���-6�'�����t 
<�_��QJ=@�T��7�ܘ� (���Q��əB��Hy�ֻ"f�A?��ӿ�\���H��.(��8�����f��A���sn�t��3���N�^��&�e�*=Y��[��X;;ǉ]�"[����4e�x\�)�Vg �)[�sg�>�h�T=JzFǚ�����B��Z���l��ٳ72u�
w�&��z`����x�� �
`{�Z�J����R8�l;���8�ׁ������{ƈ�1YT�wWP�Z2��݌̵�⦘.��x�l5k=���!��ڹA���Wr��j}�f6Z:'���+���]�G���2wZǾ�Q�r���A�5.�����.n�-�8������ivj�F�qS.> �b�7^�j�Pѱ�iI�ff���=�F���*���h��7y.A9C�7�&�@��j���߱�����ۦ\<�8_��Q�=��_�1M�"���P2�(x�|��z�I����N�p>�;3[�:�� ��ZA��vj �b�bZ5t��Q�&o����a�����dN��x)h����m�������]����)]�u��c?&����O���d%M�c�f�.A�I�S�]FF�����qc>��7b�~���N�S��g���oow��	ER�c�k���Js���W�N�Σ$��s� +�W���F�Rd�mF��b۠�oG�bd��n�{ ������H6��5s<�N㉛*:s+;m�"���T����
�B��ټ�vt}���d��k��!�ܛ�O��r{���ԧO*�bB~��T�&�����H���7W��:$����c���JQY �Tl���`s�Zb�|F�.ב ���<I�g(/��L��rK�d��|���������O���3�[����A�P2DlI�7^�}�w��|�%�oF/�|]r�2���������<���|��鸲q�Ȋ��A�(�z���V�j��{o>�&�!�]�[�TG\���n5��_�݉%�'���io|g��RO�޷�Ԓ��`�X��j��:��oTX\�.S���Bjۨ	�	BL�j��[?)2��c���d�
^lc9�}����<C[[Y�<
��Ċ�>�ǵ\n�ƥ�ć�A��R��� ԑ���%d���2�s�+�Y����Z
5��D@���ߪcgVN@��m�DE�����{�#����9�(���P�B'������L�_'�����;Z%u�h~V��hD�k�W�]�v���{}��V��k?�6�4�SA~�=ǭ��ʇ*����a��>��s�ON�RI�e��B�Չ��7��
�&q�5-�#�R=�{N��9�M$�e)��s"4|=��Px@�P�Ht�e��[1��}L��W�g�X���tfs^0�DR�� �U�;��й����RE=v�+���52��>��>���Z`�!���s""�������ɮ����D�dt� �b�&����Emu5���D�H��3� �c�1BJ쮢�>�� M���#0��B0���jS<q�ľRܯIj~7��|�`{m��5����0
���"k��M>N��]�.-��K�ayC�8��q����9yz���Ĕ�����I�[u��V+v;Ƈ\ӂh�%��d^CZ%�Ei����'���fenZ\qCO�(�6o~Y���~~a@���{6��rp��)���ܜ ��9k���2��E��W��j_Om8T#�ϪzBWl� &@��mp(�AQJ��C.�!�+Lxx����%8Ƴ�+ble4�i�~��ӵ�BٽR�.1�o^ȿH['X��_�}�f����������hŴ���O��,~Wu S�b�'��lfL��Q\`�\��\�ߚ�������г�`�[?v��j�J�����	�gݲ��-���S��v�T��)�V{����Ģ�uG7�#�����,z�Y��&XdxBR��s��<{�>
�{1�k'!�G.�qZ��]O%�����̊�k�@����s�^ ���o]?��Kk봽c��n��Xhq�@�>,���=�{��і�7_:րa����7VI��Nbk�J��gk&�ǣ�Mpϔ���|�C��L}#��j�I:�����zT��g^��m|y{�F��=^�A(�N9H����z���y/U(�^Z�t�(��?��or�ԉ�ͩU�{q�d?��]
�/&�S���bZ��m(n_�	�hOI_�-�*ߚLW��I��b@X2��?>�݄�/M�k΋����[�<J[c��8�DL�����l����������ח�_FR�I[��~���F,�c�@�n��_��j���><�]d�%�N�4aTݴuP:/6��;��hO�d�f3��@�,�Ewb��T.Жx�:9jr�"�_zx��1�N�Pm��vb@T��跻oy+�b�Lb�B;τx�^4�*�f)G����w&��C1�����=��3�.M!�}���g��{M��jv��I������������DI&����M�:���1��V�B�/�����,�]��r�^q�^��-��3����]�b��rP|e�-'~���q�MGD����տ��^�����C��e�8r�&7o�d�6ڂ�><�w�'����#3Հ>0�XV�kз�#�~�&���<�<v[�sՀ�'bU��Q��JĖ:��7ϼCXb,�x%U��V��z��=��n����9�w���ք�ߙ�3�k���Ӗ�ϏN�z@1{�b�dj��P���R|ȿ-�@I����n�5�ȎH�̩����Z���M��vh��w{�������>��0hf�M�ia��|6c�OՃ@��	��z�y�G�NL8" �{�>��\,гk�N�B
G�����p��>9R��Ǫ��cA�,ȏO��p��鶽A��.w���%����9��@ߕ�}��T�+��_
��$��jyT��+ml���}�����g��s����.[B�,G"��]�� �*� �}��#�ދ� +Ld��=���=�T(�,��肕�V�؉�}G�-?}%ӱ77Y�n��d<b&6G���911{�7lK�<��I�j�`�Y�?e�֯�:���y�����xU
�|��c�����\A.V�_��Y^˭`��E��ukl()�/����x-��6$[�4�J�,�\$u�1;F|�.�m��-�#t��6__�Πs?푅��͆��>U��\�z_׵����fe�g�)��^<������`͜�~�9�wV�>��¦UTU(\T+�k�Ep��8��Y�6��~<�ˠp6|V���	�agdM>��x��K��r�O7%D��ơ��+����]��,�x��M�p]=�e�ד�Az>��ϒ�qǝd�\���g���� &�e��Lr�X��R~��b &��
'#���B���N2��*���=�(ŭ�RK�~�B?��!�f��kW��{m��W'�$0�tK�d�%����!��o\�\�	�d�n��.�ݹ��
����2WVޞ/�"��KA�|[5y6m���ȿ~ ��Zh��q�,�^^w�!a���K$G�������4=V�7��R���Պ���ܣ�&�>)���%�s�c����!����)y�1S���+�#�띁[�7u�7�>�?��z6=�T��{j:�</h�HV����2��ˬoOh,h��\:����H��{]h�-�h�Y{�hz��pC��h�ե���k�O��m����s5ϭ��wg	�y���ڎ�[D3�eWV��ߞ�K5��}�k
��j�C�p:w��4����̬�.��4r��G_Ҕ�s4���qq^d*�4r	�t�g��ÁFB�$��!��������\����(�v��Mlm���=[�c����R��==���F�J~�[���o*�f�, U��d����F�"��n�h^���lr�����|��@�R,���߉�R�}M�>=5ސ�u9��.*��j��㤺�ҟ#n��ڹ�f��j�����5yXwD�j�vW��1bn������7O����^�q9U�Q�2�������������ܭ�O�{�&���;�ɤVQY���Dںi+�PV1 �""  �;&���®44� "H'� �(�BRBGj %y'b�?�����᜜�9�=3�~]3�=S�nk~m�a�������'d���N+�7�
s޲G?����q�iy�z=eTk9�Ɓ�6ϔh�֬��W��Q�7���P����	�o��h�x�X�o"�(T5�O)����9@��k�Mk)�xJm,�\�zg�)�
�|�:�a�w"}渼�{_o��b��(���k���� �s�B�T:��,�i6X`��EֺRT��5_���h%���׮�%�;:e�)����E�kJ
~�П|-%���eh�x�S=�3�� �L\�;�i�����G{�Q���W�y�`@�?g8�}Ʌ�xjQ>!5�B�Q�ń�"_
?g���g�G�YD��j�ܰ�w^w9�� A�å���R;� ��9���%�g�&_��}o���j���#���0�u
���~�mVr��i���4}�c��-c�o|����J;��#��A��1y.O7�2�yN�,�E��qGiU3�[3�,�k#��w6mi�f���������QE٣��tSg���P^:ϣY�m;����ч�Ҳ;d�LA�=�����D�"��щ=D�yQR���ov��M�\��-�:����i���S���;����먣1T+�k���Ç;(k�Q�ON1F��?���h���k�N��ų��FcVxt��vvxtG'���?H�{���
�6���.�~n2�OR&�Ϭ��
�6�D	��6LN�*����q�#p:Mq�meȑ�W��uB����].�o���!�:]G����Սw��='j������h'k����Q�h�Z�W�4�i���F��A�p��qݞ������6rl1��Ν�O|����I���Ɓ�qN~o���+����u�3\a�bA�]*�fα��J�/��:�E�(�ZոY'�|��%��J;C� �*���,������z�Enw�jG�kcK�����c��Ⴛ�{&Io���l�Հ�\IV	���Z�n��.����_q�V�Ї[��h�`(�}c�=�;k�j�ӄ\;+p�%��@=R��GlUMp	����Z��P~��숅4�H�~��	&�䳂N^yg���Wx%��,Z� �M��� *�%���~6�^8��h��&�\�U=Ř�hh����l�؊�z7��k�*��L_�(©v3�(��b���}[�gy��@�tL:��*�q�m�Q�qޤ�ϣ�Z��뺣�@J/[�݊v`v���ޅ�t��;R��=I������G�CG�5W�ś����gm�r�-�3���՗��t`Y+���Ѭ�����-y���vp�6��۬nk:D�)xMVaܯ��J)��U���퇂�Z�,��Y�AnW�[B�,no��2�w��J���+~V��W�	
�.�|zH�O-s&)��:�P�v�����OU��+&7�������]r��p�C��,(odh9���bc��3� _=I�$)�J�	������O�޳qG�EN��:tj�zv��z��6�n�}�qnE��y���W�8���l���U��w�*�_�	�U�!vظ%�7 a��q�Yă�MC����Ϯ�>�� ��O�uɨ?'NZ}b�4UY� ����x���ϩ�Ӆ97��R�)�k�vwu���,�>:����9���!-*�N�²P����lJ��d��z�d��\��b9ܹ)�*U�/s�Qj~h�_4�_C�r��(�YǄ��˄}�6O̒����p�A�(��,0�����t���p���Ҧ��P�����j���iѪ,{k�Qĝ��;�S�tXwwoq!�X��P���b�;MW}.�%C8��.X���z'�l�ư�5��*����be8��]Ǵ��G�;eO{DQ*q�e�-�v\[f��QC���}}�k	;0ީo�Qi�
�F|�w�Ptڄ�tz������*�}�W)S�}��W/G�T��#�yH�׮�i��AOL�o��~T~�gx�s��=�BEg�?ە�q����:��p�ۈ�r�5*(��L�h���OtՇ~'LS��=M�>�L7���k������4��sK�)p#3����ƚiڮ���f�n�y�S4싺��Ρ���JV���7�o�d�A5p<#_ƛ�M4��&��<p����*C�.B/���a��w��+��&΅eK����i��m<s{�?퐙��z�8����x�d!4��ƒ�Z���|$m���΄��2��C����/c����X�'����w0����_R�ЕU��Y�c�s��:�D�j��IAe�+��9C|�p+�G��:�K3��6�vΐ�-u2>�3z���p{ΖD��$5u��վ�G�������ֳ�v�A��i�P;&�C��G6{@�y��5J��H��O�z�yIk���^V�F�Yk�2;[�Ń�o��Q�O��5�����Ԟ�����=�0Zif߹La[��y��V���zeviK�-��	X�U�x]�N^/�X�Shk�2*����[�VzͲ�������u����u��A��1��j���p�;I��]��o��9Zխh:Q���o}��[��}!G��K��H�J�x�H�#��9�,oZH�^�n�lT�	���O���Q1�UwF��ӵ�|;'�:����P!:����3���������o�������E�����.E��n��V�\W#H��a�die�E(x�/OEsZWyP��_��V�����h����GxŖ"�K��3��K��νQ&p[t�n�:d�r	�<-�샒@���-/���X��$X��[0MN	w	TP�,�� /I]�����_�K�E$�e��6ho#������d��H�B�Z^��}�S�w��X5�MNc�y#�[l"���M4����!�4ke�s��F*Y&��`ڸ@짢�GB|D�܎Hf�j�oٸē��2�DF΅�:9v���7�Y�����YH1� ���>�L�e����9�yZc��h���W^�6�Z����1+)� Q�~r?�o�>g� l2�4]g}���O��XH�oɁo��h�}�������O���VŎ�7�,�!�QK�����Z`Q&!m^�jj��	�ݽ�@
���ҋDӡD��{n���U�XY\!��ooDx�R�̛��Nz[
� ����3�G�ݜ!Ij]��;�!�Ү7j��q� 3�dN�֟%�	�)m}^�cU�"�z�����X�!��=֞z�,*��#����6�&\я�/�p<Q�ӒI�g),�����a�8�n��'����%�k�c'���\�z���Z� �����ڽ��ўE��*�&�Us�M�"���@�6*�A�U��hf/��h2���H/�~^�W�J�����\�g�Gz�*^sd9j����@���c��vnm���ڄ�cy��2l�J(bx��xs����ݬ5�cJyOjb�'�Wt���;P�`�H���>�� t ��nX�� ��+�)��_i���C=|��`Gv`ye��aS�����Sʽ��i�Ԋh��߾�sO�x�$��T@
1;���N��ng�zt��R���(Gۘ^�%�.B�D�J�_{��cX��;W��6�6�_�8>L��7b�ʃ�����
�B�x��rf_�	�fY�{�D��M����7{�]רA��1��L_^���/t��Onm����b�����N��8�(�J
�3���Exl��B�7ǌKWi-���OH��#W?�i���	�������l�P�ϋ-E�� �W�G<$uIn������$)�V6V{c�s*��s��e��הԺ���Z[q��\3/��Jj�%R�^�;У|;0��ON����%���`�c��"O��`<�Ch�Sj��\�p�SuG�)0K�n����Os��2�
8[d}ۓ��4 xu��jB�u��?o�vR��!�}.��m+�;�������Z0������qV	#��F���C���������HT�)05��0�gP�o���G*�5���Fr�����[c:�'Sj&�Z�/����=��jjK��a�&�3����O���1�;t�m�&���~D�Ȉ����� ����S� |#I0�5���w��5���x���MoX���U���h�k`:��EZ��js�����b~��?��m��Z
M��.�x����T P��ҡ�K~�S+�)�S�W=n���>�I�-����z�<��3M����Ќ�N�bs/�a��F��DԞ�D:v
�ݙ��_Pj�(5$��ϊb���4Cn�w���$<^��aH��JOO�I�V��óGGg���%��Z�:�t�Y���df&�Q���������uʓ��c�3��q�%mɪ�;w�v�:��9 z}�-���΢���Y�U,_DJ��u�? :�~��>D��`��=�a���@_v~����ū̢')yC�����w���T7�~�B6u;�ϖF�����jVm)�Rb����}�X�5� ���բ���R�;.�ǆt��ۂ�2��_�*�3�yZ�/Mp��P�_�D�؏����3 �1)؛���,�EBV��`�ַ�Тgm�Ċ�l65� SZH]�?Օ�PB��.��0�ְ��8��͵M&T�5�3��n�����
;��&q�����0�P��W��������� a޳L4��%-�J�JmC��)P��z�	�gi/�4/�z�=�!������|Y3�:lQ��t��l(��tH�[HF1����@
�*�ݠ�L}.��-❞�d����(�;�ޥO(��M$`,LĹ�
�~`gu�Hi����ö����O��;�^�p�^v�t�1��yx�U~���C=��ʆV����i�:&�@�!o\�V�k`�"�7�Q�Z	��d��|����۾���AYW��	����h��������D�-'�f~�p�u´	s�S��N2s�%$�w�����X/���X׆�~�n�s����^����"���7�/
�'5Ҍ�.G�E/_9bϫoBV^�'����I����-8�Xr=O��#�Pm��/3ܧ�W��:�R�V�ρ��NG�Z6�<Ζz����8�,��ձ�U|��"`�)υ���;ۙa�ZMakaǾ��=n�ɪ� ��Z�7�8�������(̓_���5i5����ҹ(�|9�i6���{�}y"J^&��py ����V���Adq�|�d�.�Q;��d+����e������!�t���H�^��F��>(�	��j�J1�h=`.g�������R�?���m4_�����)��� jl�cc�G�\Z��b�\]u0c��<�4h���# �+E8jͅ�Sb���7��4*z�eY@\��	�G:�#��.<#�cl�	��M��&VƑ�Uy�y3T��h滬���,x�rN9��q��M�@P*?�%���� �ۍ�Y�:vK��.�WΈ6���t��ȾV�4Zi��q=�~;=�T��U� �&��. �ݼ���h�:��<�-������B�$�VA��{��O˦$`��B�E�b��t�!|����Fs�<Π�j�IP��$��t"h��,3��]R���zR�
�J;�{�� �
�H/|�6QT=�4��g���*�X�)(j��vк�5��_��lv���ϕ����4�N}�����k���=�n���dI�[gI��ɼ�M��|�����<�|�<�
1T5q��Bf<��`��~YYdd�ENWt�C$�����w ��*��=V�	Aþ�7����f��d���yo�r1�=%�]���|�P��h�ڛ֭�ւJK�	/t�\�~w��e����d1R�n�O�S�p�����'���Ct+�����U�g$h2�U��b��kd���n�9��hpޥ'ό��א6�� �LR���E��}��s� ̒�6���u�vm:E����-�wI_���|L�$�9wഁ�g	��H��J?�T��{�#� ^j���	܍$~��l�8%���'����b����If�W��l/J����_��TI6�.��ut1�ÙJ�QP@��ۓ��i�y�+�C��)�o�~v4_x��Vg��A�/)�������A�mC�����Aͥ�e+��'_���훊��ok�F����mҶ�DXx�+��C�;�hq�U��K@�1���k�I28��l�'���@�� �˱o����W�\�g�_���(�p��U%�����eNFi!d-�d�E���[��](����t[���׷pFQJ�#�н���R�"�?�{�B){�iɶ����+;��P���`}�`��sv �x祯Y^2clI���x��\J�E�9e���Hį��������� 0���_l^h��<�k���0b�@�劗�pב��蒪w����yF4�vOcN&un1VC�[5L����E�b�p�=��X
�߷�w�W�ީ8�ٲ�v�֢gdm[U��@(������@�Hb�e��%�>������
�Ojc$RbC-�L�;\���t�v2Ö�o����`Bd$����Y��w�nDV|v'�3��1����$ՙ�������F6񲴒�k���:b7f\m|~�$~C�	��'��v�`�p�pri��x���![��+�+g6�,i~�v`�lZ$_�>GId�SRӥ������xA�#�jNJnl$�a��pF]x��-E�jn�Y	5��X�����U��,����+@��v]Y���(Ls��p�B�`���5�s��ۃl�o����������kk}�j��|�\3G� ?$<?��ߔ�ܣ�yv7�t�)�㱏���g`2o|̸�]����5��*��:�%�_"9߭(`�A#�{h�J��?@scƾ��U�}�ܞA���,��s2Y� %(	��%��`aY�ŵ�T�����||���@y���TCW Pq\]�w�)��c��Fk�=�cU���S����k���5����zۦb̅��
�9	��c�HTG��B���Н�*u`�9	uy<Ց?���'�^J����R㴎J�`0Q�d�a�
:�R
����AC.SO����\�ꐮ��';_-����u�۱��Tت���2����;����f��;]*�8P�a���=�̡�p���S�0�c�g��KqթJG���d�!<v��/=P0��w�^��-�qxd��+,J��=�@�eg~��������c�����:х� ;�񷶋�������U��7/t�e=��AGE�����Z��٣���a�k��;ZU2Зt��@76�jX�����XێQ3ŘdU��<��z��@Sy�
`%lӗi�<��V��R܀1��&���l���K�
9���h�ip8:%f�	�a�3������t�^eǳ�>�7uԠ���9�7D�ժ^֎���c�F��k��!��}8@�_����:�4jҟ�#�M�X��g�� |G&C�}x���3i��2~(|Z�<}���@�T�Ԯ�MW-
'�j39�B�(M�d���rF������`�����*���?�y�v���Tɟdf,Ҿ�%PM/2����WX�����?���F
"3�D�Fn�ꇻI�vy`�o�v�KT��9��t9��Z���}�O�k/8�x�y���V��B&;��m�QB���T;��/�������8�F����+��j_��ɷq�։��&>㭝�P��(�ϊD��Ξj`��f�U����g���˃ �R_|�B��gYi�n�d�)�߱�m�&�Fwڻ}���&]*u�H�i�@Uw ����mDАzfE�^ h�7?}PF�v�����r�^;���͠���Ϟ�*[��N��	{wU啨�k�)#��c�y��<븀�[Pġ���*�1��	N��0�]��m9�ۦ�i>v���1�M@`h���ɷ����š�����:�����
�9`���	O�b�O�#��T�+]���X�ۣw�|o�����PM n��������`�%�%`�վ.��$ե��k��?�LXX�X��I|D��|R��h~�C��3�����m����g��9�A�_l�+�>y
k7�[
�~_z9�R�[0�41���k�������/���;�8ɷ�gէ�(�j) a������b�3��9��!~?��ޞ�yH�_uW�m~M�m�dĝP�w��@A߉�q�0�ThՇJ�R6�0i�]����ݸ���)�v�Q�7D [���#b7��x�䎈�����u�]0�*V�{���yA��l��jAo�l���M���.���y{PUӎ����cƣ��ɌۣyS/!\�۱��+��	C��]J)�n�z��C�+�綃�4U�P(���0ӺB��кݤ��;�ik��}���U?���/�1� RT��t�B<�4;�%���Qq��R�V�Bi/l�?���{-Rt���&�~����/Fo�������b��9�߭�o��w�2>�O��I�2̹���?t_�_�����l���u�J"�%Pj����c��N��T↲��'�a6�:�~�7�U�V�ps�G����|��
�P�\X�JѤ��ٶ5�����(�D.�Ү��Ry�/X����b�n�$ZR��6hl������U�rՆY�0��Ü��~�t�/R���s���,�ٰ��I�m��@WYت�:������S���꠹��	s�;�pM�J%�*n���P9��`�b�~�n�oǋ���^䭀�HXз� ��*'�A�z9�DK�r�>�n�+'^κ����M�!��Z�X����*���Z���Lت�Z���9)�|���=�ɝL:�mK�=�*�����F��5��~��[���8�4�cV*�9�Pp���U0�z����_�L0�c�O�tYD�/'{�����mQJߋ�]��5�O�VuHf_T���+���L�9(Ka�a;���~�aJ�. �L�!�1=!�.jk�R)s�դ���:X!,H!�>�%�1��G���ErT��i*=���V���]��cէ3���~�������+��u�J܍�oR�?���)��ѻ�{������=��G������n�R�Z�5��uw��'�����{����_�v]����K�9���K�U��~�[WVeo�p��kW
���~Zxy/���R�8���K$$���i�b-��I\L�X�HQ��YI�M�֣�"�����u��߷�Y��ʲ�\�����_������&��}���_w��o����ܠoj�b������7���ߠ���{��|��0=+Sp� [C�,��Y�e�X��aج�J���p�t��Џ�+H��!b�?>ν+����ܘl�1��m���'l��g�k�jm�7D��!	��#�^�'���v�����XG���<�AF�nkv�k��3����;?�8Pi�p
_ٱ����$���H��3�H��;�%�� �9�a[���y�'X�c���UXD�Џ�W�f����o�^V��hY��Ս��^c��G����O�k���y��T;�$#� k������"J��@j=�u�GB=���`����ˉ0Mz_dM�ZO�@g����0���0��.�}.��iz<H�C����������+T.�}7�_Vd~����>���Љ0/�`)�j�Stp�#�\���U�Ŀ�t�
��Vy�Yi-ֶ?��!�o���׸����ūZB�)��K-ўG��M��\ޮ��hJ��k���wU�\EV�@�7{�K���pw���E�k'����dԍџ���/
�z�r�Fk�\0��.��zGB8%� ,��Ǔ�Ex��������KE�q|&L"V��R���Ȫ���:b>9��%�R+`�|#�/��1(���\����ߠ�W��ޤ�2�j-Y}_K��};)6�%A����ydU��H�0Mϗ���upCtZ�U��,�#I,���{丘��/#�r孃y��������cIC�{W�Md���ȬC�e�Ø�O��ǹs��x��/�O��~W��Ӽ}it�r�0��|I|��S���B��_�I������6�:����LDz��h�2�j���5�x��q�=��ְ����J��Vv��V��B�Y�Y����ar&
����y�A�0������gFڃXq�zkJ��Ү��+=��=u8�S����z�:�S�a8~�2o���j(n��,�i���D��߭�*+�B�&ۉz.n�����D���S��u�fy�u�t�~�/V�A�O����w<��C��Яϡ���d9�x�=Z-���ch]TgS�/H������%��F���?sN��׏�J�ԥe�H�9bS�۽T��Q���0C�h�}�'-��6�._�~�5Ab�ǽ�.�4�!����;�����5#8�|�<�
ѹ@���F]�ΦK@	����� ����{�@�D�����\�_�^� 
ٞ�����~s��T�732����&4fh��f�H�F��j��&E���K$�#����`p��&e
&e�Ts33.0��F��#_#��z��܌x���㹧�4?/Q�¨ "lޖu�X|�vM���D%�����hl���w��F����B�G�Bm�x�AIy#њ �?��F�������ht�W��!�y*D� ��Q��׭,~��b�H��չ��XEy�c����� ��O�|\|�̘��C��m�=��-��}5�_�/�f�O��9ЙщJ(ͨz��v͎�H�,�L�eL^R>5�uZ@�Ãl!�9�G��N�Ώ��mOG`^:�-*T����jk��4��eZklL�=U�O�ℬ�纭*�z��2V2kr��ҽ'��
�����f���z�`n��ג������v���	�"N�w���$���t��QG��m�W����l&�3�X�#U�	��4��ҳשa=��	vב�(���IH��x��N�I������e��Z��'�����0��H����K��G�%]�~�sw���5&m��2����'X�E
�軋��6���IGˇ֎�oyq)��t&6��D���)�7�*�gG*��_�����B͵��ƃ&5}�g���O-�Qr�C�C�9~[�^o���!uV�}ɨz9SP�~�Q���.�EƌT��j�>�t[!�zN��^&��>���;� r&��Q�?����}���;�n�NSTWj�6�YP^YT.=e�j���v�O�����ƽ��Qܪ=��p�X�o,f3�<���Ks�{��zY���&K%OR����T�kF|ԅ�6��M>?y�s=����;W<?~�-[m��B�N-��������e�wTh76D:3�dٛ���㘂f�r��=9���x�����0�����\7�e;����$����-y�ٛ�p���|+�Z{Z�0�X��yf�3$hW���A�|(|៾�Ŝ�`��Ǐ���=G���N3�~r������=Fp}��ږ6�5��~�o�~�޸"	���˪܏arDS�/�w��׭�{�4\h�o-����4SA�������љ�`C}�u/?Q��	u����ƶ���m`��j�w=aaa1Ӷes5�̱��1�Uv&vw(u�G˃!)V�>�6um��;�2U$��]a����'�iCް�td-N�t�����b�G�c���CD��S:K�b,����¦H�&vh�|^�x�6CJ��03���I������3�0��"p�KPbl�i�A˝�/����;�,���>Rm����7}�� !�N ���Š�&b
�o�V��0���B�.U/|��jk�j�1
7��6
aA+�8��s�v���N>��VJ�v�N�{�%m��=ruv؀u+�~|AD��ԫ��Z�Ǐ�>��_�t��z����uX�Tz��փwiʵ\��̣Ǿ,k��OH�:�<W��p��������#o�;f᝸O<�[�v���ȸ����yI�nQ���l��ϫ���t�(����(1��?�0��a��،0�&���7�4�X���;��'��
Y���u����6�m�M���1��-�{�^/Ƭ����GH�[E�9;��͘���G�S�W��E�lǪ4�h�X��P��ŕU�VL�����b����f16fHq?�w��6��sni:��u��ü+�%��̐���=�d��{��� �*�pD�}���Ƽ�P·c�k��;n�1(�: ��֑f�6����ӈ�f��Ѣ�"��x�y#��M�c�Ew���'�L��x�#a�J��o� y|,Xn�����ɆtƑYEI|+Q,����-��c���T=��i21��) �h�-j���];�3sV�Z}}��̈́e��6�
�sUj��g)�v��g�� ���c�����)���'*Z�&���xX�d�m��-^�(
���{W�˞�����&P�E_8y��i]Ů�7�� ��^q��`��7g�t����E����:���&Î~�&N�b�ոR�r��H>�qh�7�!g���͍qێ{Ot|E0a"<���qz�k�٭���"��7HD%=��S{A��&V�x<<"6��A�D*l�9}$��2Itt{���[-ڶu)-h��xI�ܔb���t6�������y[�~�uW������U:��p�A�K����/II@���J�bٍwwAw�g�Җ�ul�u}[Fr��c�vr��D�G"Q��Se��V$ݓ�v�/�Q���֩Ү6ƭ�Fh+�����_fؑ����:Z.|��CsGc���.��W���D��:��w +�1�m���T�Q	߫͠<��+�i:���h(��T�]ʲs.�'��(o���A�60ɜ��ı�����r
��~��J���b�����b�ѥz�N�_�@�jܿ}�x���^�����iْ�s�/���N@�9���j���9;�k]�B�� �u�h���"i
����7+2�qNd�M��;���:8���<�.��jv�h
W�l�֭w�e�ΞSk���e���J0����b
�lD��SG.�R)�˙���!�.��������g|���Z�PQ��_nY�𳘟Zm�p�Y|�3[m83M�������l�v���6�������Y���W��M������H���������ƩI ���������}���k��ǳ#˱����u&�,m��"����/=5e��C��&��8�bE�}m��Sl�7|�*-R��$�z��31¯�=®H�沞��[Eix��4�bfr�ֲ�@e7'�Pl�1<w2����n �/r�T-S ܱ�'�5�+bC*dff��n��l�����6_	1#[7/Z���2��l�uFk��7�R�HR<z6�|֐��.��m��}:u�j'��q���˟{��*y2�(6`e��+���j����TH#�⒎Ss6��s�/��q�r	��A4#�v��xeh�MZ�CD��k��4����T#U����fUb�*0`0r��B�ɉ�7�H���X$��-�7�^&���ނ�˯t���7����T��sEw�����z�3��BCZ2��9�l��0���zO�����ƊTؕ���·�Ӧ>pE�O�3�(��?��H��(������Ga�z��`�:�S��O2X�Jէ��� �� �� FEE�x�޵��Z��T�p�T�k�~��N�r�ƋD����l�R]A���v�����El�٪��Eg��e<N�Iq###^�VhM@�k<z-�M�������<u0l�Q�<}/գVs"Q����m�#��u�L)�̄��6��դ0�d�lh����I�]�iW,�jΌZ��`Yf�DW@��pC���q��K���ؗV�~8[�<'��֌��(����l�x�x�������3����#���J�j�0���NO̎�F9\�bdd�{,��k�_��@&���2b��B�'6�pjM~����!�ĭYq�!؉����f���vu��͆<�X�u���3�)�l� ��m;��V��-��b0�\�K1�lg�V@��>�Z�"�^-��c��(`�&Y=���t�?�4��y����g��m��		au��'�e����C��8Dw��Y�aH(,M���)��F��'���D�#E{vt��O��d���G�*rީ�B�ϳE��B=�����М��G������.��;s�|��v
'�ΓM���d�z)�VܛQ�n�.2P��ܺzBfh�du1�$��[r��zT�P�h�B����y�wIG�Ei�wb�{��KW3��C��m��ز�q��3���ͭ����k��d�����v�+qAeT�8���R���xc���5�F�֥O���GR}\��r���8=�ˌ�?���_�Ƚ�a����w�Oy�+
\J��ZY�3۽�;X��X�(��2��&N?4ᭃ�����Nd�R�����ɕ� m��G2PN7wb.,p�f��G�&5�8�mHSB���Î���7n̎��-�4�P����x;I���6e2"��^�cG׉�Ӧ��_E��H����$G�d�x���[l��a�]��wXg��B� �Ϣ��r�Q��˿z�x��ʹ��9C�ɕ�
q�����0�Q,������نS,�,�[�YN2�4Ҭ{e��I,8[��0�Z�j&�1���:��Hp��7��uk@	kR;}8��'/�H�k�~+�0�#��W�?� !s�x99y�ρ�bG���hՃ�ǋt��3q�3�^.ڣڷfgE+Z3��I1���&Dg�Hl1s5�z�Ԋ�!&��ĺ ?v��&.���yj/�&���!�z��w��䩦��*:���Tk�R�h�(s���c��Rن ���g#��Ht�I`��:�KP�B�H���de�a}|B�AT��ȡl��<57*?�>ҫ�1�𵯸wW��>�@�s�*5`H)6Xx�X�6Z����'����!P�X�}b���U갫�"�=gӈ}��E�~.r���N[�:[�}�1�,"���RV�.�"+A�&Kž�W �`o��|;��]����.�)+���%
ss-0���1�u�,�;^�R��r��3gj�w���,\��t������ u��l�rlG���\��k5t�h����g�N7����u�/ӵ�'G��>A�8��}��n_�)��Z�>�1e�� <0��[��  <�����z���ZZ�����֭���<�r����v�dk��j�����K4�� (<>l��^Gm��LYz½�dz˖|�S�R�ԱH{y0�R�o����J�>ޮ��w��U���%�Fk.j��yJoɦ>��_LrF��73���V&�dm�S �����#�����_{�K-�a/'�^_#�������c)o_�\.���&6i]1�S��oO���n:�l������Hi�;L>�Zy��Y߹]gz�C�i3b��]xP��O�$5'��&v���IDr�c��,�����0"����bT`�;���9u�P�����#yt:��z��R$�lD�֝���F�HŨ�_G��'���t7[�ZХ�2��J|���6�1:��|Z�{�@���G�D�߁��E�ϒ�:U@�ḧ�z�<�8�!lc�����Vd�G�� r���g�XZ,dS�
���y�x`��O���+C�FN�����jWt�n��1S����M z��?TH�y>}�[?o.zL�
y^'u[����Up|��w��x�:t����/*�EؿM��P��8=�Q����@�o���Ʋ���
3xd�3����{͎}���#W�T:T��x?�J_S���h�|�f���g-�˜tu���C.����ܵ�f�Q�ٳ.�}��=s8���s��l�&{M�k��<h��*Ӳ�M�99X�2��v�N����_c#�٤���YNT���^�:r��)�XF�� �(��3�^�Dr2e��u��n9�O���D�\)$:�����-�ԩ9�Sd_�IfԄ_+��h��l~���"��CV7ӧ>J��ؒ$�x+�`*="��]��3E�w���m,⹀�A&�א{���cE^��W�Tg������Y6~W U}���w� q�asxVxߌ�L�Ԛ|}�qQ����T\}�q��`iI`iP�Vd���=�������Ҷ5FK6�5��#����4'u�Z��D��:��"g����`��������<�xw1����af�x���S'�N��>�PC�ti�,�0c�v1��D�Ym5�����F"-�&_Ů�ǹ�O�׉�lz�lZE�+�7�(:t>��w�V_��ĕyi��p9�`�)�u�]J�u�.��ڝ���h���{�6���������t��a����:k���sV�u��AG�P���>3���s�*��W��W���ڭ�V{B�,	�}��(âp�"9F�.�[�K��=e��Y�T׼d�:Ɩt/u�:�e��[b�Ѐ��^
���h�ň���
*�@��M�&'�3kD/��5ֿ���j���Td�?s���$�\�`�:���@�+}`)V�����ޚף����;���?~�����H��Wr�%?�y���Q������ ��.:kw���a7��������Q�F���SMYi[ۄ����P;��!!���6��jںty�����ӟ))�<zU����jM�A��hҀn��9.�[�}wZNY���~8� E�J�\,'���39RF��+����S�a4�$"���Au��07�#�~j-g�1/N��흟�v0UrF�m�ѕ���2Th�ӷ�.�!��7b����K���D���E��r���έL����~����k���-qb�fRY��F���n��&5����߾Ѣ<��X��jzm��)�9/��t���˼�4��O�S�h&���"E0?C����*ͣ�-]n�S�s|�y�fv;��^i�ExI��Yտ*��x�zt����L\|��� #C����yB9ᥣ+ʓ9�~��u{���8t9&hם��ԫ��6[���;~qʋ�X�����棑Lv�P�+�P!�c��_��n�{@���&_� �I��j˯���l	�Z��mU#�߱��[���m��%��^V���?���u�D)/]-�-P�'���4�Нyۈ�@%��ү�l��~���c�DC��exS�DF��.
�,��<`o�)�nU2�i5�Y���x{ɾ-_�FY�} _��XI>�S.gG�����j��j9�]�2�vo��df�����u�����%�����I-��=�Q5~�s���Q��Uy-ܫWR:!k�+Kw#��W��KW�4g
�;NNU�`�:����:�$YM]6��m��c]�*L�Yۼ�\��^�|��O��|={<�l�0�DV�>9is���I7��S�Cb�]]�`�&��f��d��_ܠ����3��;g	�3
����J�X���= IEF�
� �
�]7���?�}wTSY�.�ʌ(̌��GiJUz��`@�"ҋH�%����J�Ф�*���%��!t�K-B�;�6��{���Ǹk�ֽ��}�����99{�U�{k�.�U�%���'lX^|	���C�"f�*�񯄔[����_�bkg�ϝSQ!�)x��񘅂���2�	�,I/��-�U	S�
C�Eǀ�A��[�"C~fы�5��+R�d�G����x�Q��cH����fg��62��Y\�U8��Y���{�3�����S��"鉔�j�t=����&+���I44$Ǖř����NuX��>s��R���Z��V:���n�8�ĕ�^g�	���c�#�J	,�/oR����U��l)"��M��m�n��I[��@i��}���,����,��S������΃풄Y��=jl@�X�}���9ys�:ć����!(s���@�oْғܷe��+v~=	��h�"�$#S�Q�r�+k6c��y~�Q�T-�Y��\b�R,�1��C��K��R���]>=���$����k�8+�T�_�3��Õ�$�_|+�j�teS*#��L���L���L�[Aju��kW_L&�DR�U6��9�Qў�5N8�Ak�bO�RxK8~g����� �X��@�%��uCiW�rmĞI�-��rJv��U��/b�[yz N�^�,�֧a��R�4\)�%�,!���G�4c�F��!��fE�m-
��L�⥸�m����ع؛�d�3
yg�-7��ǧ&�����>ed��=2�|j"E*���4���{�w��y{ϥu�|A��
����ZX�Un������4�I8��v\rʑb�|`&�������#"�>G� ���*�w�q$�i�P1���c�G���Z0;�9��_:R
c��,tN�m��*�A��|[�irO9{���a�}��q��V���0f�5_�}���`�H0��&�����}C�Sk#�.b��ڜl9�A�i?5����ݼ�����Vz�l�A��4��5��C���ة�8n|o����L�bom�Z�L餄��5��؊��������2_WȾS8@k��_�g���{i:sf��3.�U��*�vU��{3�Z]J/���v"��V�{�2�Gf7�>o ���+�{!��O�I�q��OiM�NU(�6y`�������<��l�f� c���hu��O`�3��N���X
5]&׷_c[��$L�C��0W&�
~�xzYH������bs8���&E��W��6tv�2�gt|iqW�O��&b	�E%Q�ľw�9d�;�*�R����� �v��v�]��b������:㹤E�F�\�d\�)hc�B�I>�B�:�R��A3���T��k5��]�
 ?ǈ��?��7�i�1�O���h}�qF���vMXfu�f]�B�}����- s��^��TY�2{�j����l��F��^�7m"=���^q$C��1���U.�����X����ä�yŗQHW��u�����%��
�d��{:�6V�jS����읾�fmo�4��Ky���_��`�k9�E��T4�v��N3�+P�I�i����V�z!�6 %�����#�B�=xJ7������*@�ϳ�Q+U�T���*B:���Y%�Q#!�KP����9eGC�������edm��1O��ثb;�m,�����&�.U͗n��$Ò��U���i�7e�iC�:�k�A�H���d�q�W�%e~9��-(ϩ�E�+�d0iA{��ݼx����Z��c`��Rbe�	�i�v���4�V��,O]��'������A�v)0N���!~_��(�Bh� "��p���u�l���C���]Z�,����fK"r%��D2[ ���:�[B)l����/�R�I����eJa��X�*Dm �ی0C���</�W�m7��1�x�u�k��e���J�h�������0�IKF��w V�H�פNj��V��6���z}���,L���<�F!ߛȇK�(�%�m�6�jCG�XK��!��}�_���˱�V.}�'O�`hVزN.g�f�λ�	�ȿ#�f���n����s�|�7����V�@�'(��z�%�f�a�ҍ	����|/:";":��D�%8��eA�Y ��p���-I���`'�s>��`+|���ľ����g�50�IX����os�/iP�E*6�[ �ķ�9vr�o��4w{����y�i���}2�2�/�r���ϋ%�?�X��ϟ[H�%[�19���1����6o�a�"��:����M����b��^��Y���^?�cEY��y�}�a���-NVc�/<��Ƅ{`��Q��g$�ك�b�rb#H�]6wʕ*k"�J��Q��#�t�Z�
��ZgS� A���LU���IgK�0�u��P�A-�7B�/t���#�+x)�D��f�%2Bi
�}��6�?a�'jv�G���K�re_ ��>/!���t 2/e~�4,;b���,���E�:�wߟ�Xԡ:��0C��ϝz�
��״�%Rn�/��M6���7��ч�Z'�X���J��0_�t>S�݆�5�t4_��Eef��פa��G45���%��o��eIN��k�?�`��:�vAg0�1�����T��9[����:���X<OKSV`��Ӱ�7�Fs��ge�%&4"��UW�<ȣv�	�sM�|Z���<��|��_��[�=4`c�?��Z�$Gt�ض�zj˺�U♔���B�%Ӂ��Tw���R�qc%�''�b����,��V�K�+,K�%ZA؇[�6��:7�>l�ͅ��kwp���}���G./h�
/�~�QOi	)8p	<�Cά��9��չ6K���h]����x��"�?��ㄗ��gErE�m��%.>l0��nc�C�ͿҾ}#����Km� 'yb$Z�mF
Q�ăw	���(�SL�=6���^'�L�dĚݛ�ȩJU�pd���X��}����B��1� |M��D'��K=�A}0f	|��>;0'�p�����`I�H��A��?�j�Y�#
��X��0�mr�?�?�$!#I �_v�$��w��C�5���HJ�Qc�Vbс\�ت�h�K���VJ��t_��6=�ad��3@�uP��jZ�kkS��!@C����c���?J�X*s`�͂���G@�Q06d�C9��G�= r���S��G��K�J�J�Jd �S��V[�rK�5!(�0Ը�rb�@ѤT���S_]Mԁ�f5�����EqV9�o��k����r��q�CĚ����LK��,�o�ì���$u�$kv^�P�pb,ϲ:��v��me��𯀅 :Fr�(�VtT��IG��1�I��II^���~�wx�e��2�l�Td��v$�5��O�)�dǡ=�ͣ?M	��"L�m�9�O���
�|��c�~T��d�%sCα\�igR�f��] kt��|� �P7Tn [�b�.N�5=���FqbB��4�*����!�ӎ[���z���s⯿���(�\�+4P���h�]5nU�V���Z��$p�Wl��<���MԿ��&��_1��ӅBa@y%~ji0�r�X�Fx�m����hq�����复p�(���6=݊�K�O��{y��e�N�R��n�s�B0G��M:�cD>?�hEN8��Z����k����7:��%�A@�z���띰�н�s��U�<+�>r [�bܿq"��%뼅���53�!��]uD?l(�6y�l����ξ502!�'�*��\.���AG��5TV���v���]� RB���"���!\�5��K���:��	�z��Dߐ�P���*�Y�O��t>���� �t�%$�u��]�r�U�����L^\�N�'��n�I�aaH���(�&H���ף-Wqd R�F�E�g,�ۣ�g���MC~6���)�-V��F��D&խ,�T��`[!�'��ݙ2����\8�
�~b`�a�ײ@�ގQQm7zt�~���ᆌg�X����T����_�LfR�����������P�e���R?vP�$5ۀf{y�n�v����� ۯ��wN���I�	 ���p^�����g̖�bB��g9�� �� 9��!`��5$J^��l͚��2|x���^�dY:�t�=
����ιlAgT�V�I�e(��u(���/E'� ]�E�U�Ax��L���k���Y�ma��g�W�ߗ���Ev�I&^a���T����~s�쌝~f����%�ߠc'Z�"��p%ء"iP�#� '�0zYR��7�����s���j�#��
euK�J��v鼉Ѽ}
��c9���fٰ�@������r	��?F[��ْ������Nrߒ�Z�c�;]��U��	�1K�D"��I坶2c���	�2��}ƙ�$.F��HB��u&`�;�F��lՒ^��g/�w·f���D���)�!���[)���U�r��&��d���ֈ�Vt�`I
�Ꮝ��}��fL��u'���C����((lN�|= �3%��g-Rf�Q�z�{U;�!�4o��|��|�u��^|�.�q}��Mbv�ِ��-�*�x�N�C<�~(wE�~���=�t���?x㇮6�R����&v!�&6�i�+�1?�`E�dy�N���`	��G�+�F&�l�$�uV�X_Q�1!��?�Q ����tܛ�=�<5�;�1~�	=w�����9w�9��(�?٬7qП�b�����Bh���u\Ql��[��8�?+Sv�;f`с�Y����<�T��]�_mh��1J�����n�OInOo���.�8��D�� �=
�g/�{���y���	E�/r�ʇ�^��t'�'��2S�k'�w��#>K9�b�^��^ �߁8y��v��(�V�no����T�+�����2�k۱�}3���]����;�|���� C�F=nص-<xF;��'����a#Ρ�3(]7��s0�ur��������A��+)����Y����:VL�X��4�c����{�]�M���]�����c�ķߨv�00�߽���ҏ0�(��Æ)�n`�qX_X�c`�Co@7s+)�G[��g���r�h�<���Ew�+S��pU[�g���s̫�Q�j4��ys��bl�4���mA�K��H]f��8^4\b�l���Q�&�װ�`���	ҳ&V�wW����|H����M<Y6���f�� /	�5���U�L%��֌U��E���z�OZ��C�%���Iʻ�&�W�XD��T����x6��L�#�ݷ�"� >���������kh0��ſ�y�6E{�)�LKԵ�����s�������Y�'�W�7����������7�Q1�n�e3��(_X���?���x�Q��Usi:�t��ǡƫE���ǈ/�Q�"`�\��&��B+����^m�#�7J��Ubg�GǖO��
~kn[�>�\��2Wn���GGl(�WR,��2i-QG8#�hhhP��k߸{F�:Mz_���O�'�t�����]�	�ί~��u2"���B�$;<j��#��y�����u�5YQanL� }�7Hy Q��f�x�ۇX�M0��Ů�^�>��z��m1]���Bm���-)�ZqBb�����ٗ8�"u]��7����y�����7G�*:珷�ו����w��r�VX�s�Zec���O8p�@s�{��R�$���:�r���ͧ>�D&��C"�l�)[1WJ��'=$Mv9��!9��������=[�9��?������-���Q8�wI�D��>m*��Ǹј���#�h�0��
m��LN�����EK�	ԶwrlI׭�1*o�
����Sg9:�9:4J�[�+�6|���ӟ�D�1��cFz�cAԿ�J�8��I=��^ͯU�`��5��z��t���޾ҵ�PW��3]�� p�`T���*���b�?���e�U���[J�U���BD��Q�b�E%��F��T[.�%�Z#j���
���`�ɭ��ﲂ�:���%!k���i��ѽs��5c�p����0�,��t;]����3���x|Ւj��_���1�Ѡ��eV~��p�Ɯ��)H_��CҔ�+j��#�(<_S���#VM�]?6�X�	�#��^�u���N�������ג��>�Ȗ\�� `��P��C%*x�{�e�/$�~��B�a�Q�~��0e�8�x�OZ�3W�/@��X<϶3�����b{�Ў�h!�SI����K���նvC�W�ФF
��#����{#�D�;_տ��|힁��ӱ�?�����������C]%�{9�Z��H�pZ}=fM�<�E�����:�|T��\N|Z	hF��dv�bvrx�7���U������zpؚ+٥�H��>&殄�X��j97W��;3�R�[u��PU�߄�'�CI}�'�	�F����D�-� �ؙ��
�m±�I�������ѝ|.k�H����r�%K:(������k����Gn{q��ԗ�N����N�"h��FY ��2.4�$���Y�r	����;*41]c#&�_��n��&������O��A��ผ|'�O`���$9�$cBv�\�$Q���O��B�O������F�m+���fw����~|Au1Ȩ&ȯ8��0�+.Y�������7���<�B��xG�r[�=I!�*�=���^[�)윞�Q~��\m�t�k�]���{FF�nt3�~�����3֌
q��l~��r~�v�~}rL����񄆛�G_��;@M�61�
� ����Jx�/��ݰw�Ǭ'i*m��T��Ֆ��2NgP_�dө��J���-}&���`>b.Y�㱖�A?�l	�u�'�je�ZN�oDI��mϔ��r�KZ�&t��3^z;�၀��ͩp��;��F���k������q�<���a��㭯;��	���8F�kz�(�����8˭b��:��ma=h{��y<Ι�&���Z�OVI��u� ����wW����_ݣ�V�E	��%���	���b{�{}�~���0�����a</�[�:��Nd��=�R������P�+�zsS�.E�Y�����j$��]*�[C�}҈M-c3��M��SRN*F�FN	:����N�E� *�������.挪h�"�d�bG<O�_���t��d"��3㬻����@�7����L⁰���
 �:q�ph��ǍɫV��A	��")�(m�Q�G�`�>%��Í�Tӿx�(-��k�y�RJ�O�%L��a;MQ!�d�s�_�7n���.�!c#t�C��.�*���K(�0Js�R>�6R�Niŭv�?��嬥��j��iɏ�|.��~�9��]\��E���r|����p|cw3ajA,��wT_t�>�As��n����=k�DL!����,T>���M�.?��
�{\{�nV��X����d��&���I+)����I�|��
?���vbb�~Ѡ�ʤpۅ��j�i��B�2 ~�U��߈`��9e4zP3/��Z��	y ��1Jw�}^����P��W����F}����3f�22�:h�Ed[E��t���?#0@��x��B��+��Q�:c���Jo���E�Y�R�@�lJ�U�
H�}E�M��$�b�#xV54�aM���&�D�f|)�j���^��D�Yť���t�@��q#�Խ�pd�el�I^���
��:��(�3[�W�^Ν0?��ND�ٷ5������&���"@��w]���0����gE9�\�WYVh���-�P6�� �ɫ�z�QkfC�_*��)������+�{{�G��>[L���1����9F$%�rcydDp�P�������{ :f��AY�i�\�hZJ'x�:`o��.%2��7ҝ�l~��;zͨi�]uA sw.���('��2�A1��V'U�fb5�t��]��ǒ��[� �,)X�R�,����jqd���jͯ薭��?�������
1�v��ܝ�AL��c��_�H����.���t:ºwP5�tB�y\
h�M��Xd�0D| �FH{ڂ"��W8���)@�D0_Iʝ�	R��b �xmc�-�#`��/QgE-J���ө�Z6#��Q�o�'(Ջ�4��"�Ծȅ|d�L�q�0����H�~��V �Bt=�r3�(�8��k��~��﶐�,6��9x��9-T_duχ$Fv!遞�&�bwʕQ����p�4{\�~�Eww(|�`�� $� \DZ2��*!�kC�w"���,{���[�\�H����H�M����;�_ �fT=z�R'<�[�js�^�3Ŗ�N��}��:5�&���owXq��adû�ƶ��6��1n��هa.����� R�4��kVN�J�v����Ɩ�\�
l�?h�bc{(��)~�plHg��F���ܟ2��X�5��@	�� N��F��"Z�dqt�B�_rCƢ� !���&/��
|k�r���m��wf�KB�8��W��4Vr���dw��,��ꄾ_�as3
���I��6$��=V3%|������Q;2~ҟ��}�	mS�5ݮ���<�G����~X��}���X���������z��˾¤��;%�,`l��D]�y�e$q�ju�a�-�{%B��[;J'�|��-OtJ���o&̨���N;��} ���>�CDP%�pt��K��}F�`Ji�����:�8�E�*����W8�ݾon���|e�6��z����'!H"3+�xC�:gC�Z�����ݘ�b�UT�$�!���=M!�&�0� ��Bv���P���u*�8)�vF��5���oWq)�GF��yĞ;C��+�!�H�+�$�}[�I��J�s O��*��»#<s�+���^-'�lW���d��J�.aT��B~:`��lZ�R�@N��.���|�q���Ҏ�^X�����Xo~-�~����<����������s���K���50<G��ߓ���13�܉q&��롶>|�E�@A�1Ζ��gBˢf�e%O �%���w��i���˲8l��!m�vx�M7oT&���]/꼺A�|2��B
���ϭsԯ%�����d�}é\��&�|���@*��z���r6wt�4p���w�N�\4��l�t*�Y�%l��.}PA�\�
MQ7�EEq�<�WH���B���,S��o�qE��!��-t�nݚ5H�.��;Й��M�8]����@�QQ'D��C�I��SF���/�&��^I��U��$�D�	��P\!��=��,����ُ�hV�����	W/�}3�&�ݺ�~��@���%`D>G�sT��1��J�l��������Vz67�r[�8�����i�=�3ޠ�h�Q7��G��Nv|���	�B��g^18��,p'��(�ajK,�����$'=̊���.�V@t�b��^d�\?�󴈝�Ln?n �Fk�r�r��nږ)�Ai&XX+=ۋ_b��}C�>���N�����( Z��x!�����<Q�Ņ���.(<���;}�V��X1ӧ�4.�\�<��V�0"�3P�d�ZN���Qͅ��&=���R��.�j�%MH�A���k��t����/�&T+'��t���:y�<���q�d	�h�ZG��I&�ؐ��uE#՜A�|_6jO����tL�	7��Q-C_J,t(l ��f��XY���C�b6{�g��R>ν>ś8���	#r�:���~1fl�()�6���3GE�f�ៗ:/8dgr�D��,]~�=0���/�~^Ni:?���U���^�2@>h�b\�
��J@1���v�����E�0揾'��܇|�,�z���bY
�-g�GI���� [��k4�����]�5��+�J���6�f�ʭ��8�PA�m��G���U�r�Q3�x�hذ��0�c;�Ґ�T"�+@�k{�~���-��,�t�����N��������__�δ>b�*'X"#�UbM
z|}��]>�����:�nL������2;	�ܫg�DlyX��� ��Q�{�'�Qc�!�Fh3����g��*A��� �1T�5�K�vQ.�`^i'n[������M����C�W��E��8�蠥��&D՜�Y��j�t���=��~`�Gi7P)܌�kM	�3����Z�6p�����~`�@�F��X��L���|���܀e�f\�o|g�\٘��?����N�Y8ƍ����/�T���($�0s�c�UÔ��rCB�A�I3a�'J����f,C�2�=W�X��9�����A,v�k�J�XQ'�jS�R�� ���g���ܺ�N�*u��N�����N�]>BI����W�N���}Ba��y�6���i[�~܁��E����tK���?q�Q�/-o�L޾��I�y�Ap�$���!~Pu�cD��q��|��Z�AUV��,Kl?"s�匧Ⱦ󏩾�� ��R��U*���X����<��m��a��95��O��uބ����#�-b���xG��%�l�"�fuLz����eַ�����#�6-R9��Т�=���_|�@�%����N�u��َ"�����N74�������S?�g쿌{-��RK��@�B�7��-�RlK��j�J�z�	%�ͅT�H����|n���O�[u�%��]����RF����k	���}��=��`�g�-0D9��0�x�������5��������!�֟rK���%�(mՋ#���i��o\��8|���.<3����o�"��R�$QQ��rG��ϻ�������C��.=��1���9 �tx{���̼�|Ҡ���'����ڈ
�[����b��yC��{������0��q��g����{��������=�?���:̊���Y��M�����jǪ5��Y70�*��;�p>�$3��Ώ���uF:yƇr}�P���<>�
���9�EBp���<�]O�
?>J�b�s ��&�Dѡ�g�4
T{S���QS���R��|dj@��b�@�4���t�p�y�l�/�Q���H�\��o|��}�	�MM��¿5<�t��4��:>)���É�r/�e9��?�p��r��������4���i{�r7����Q/�����2�K�k��7�"�0��`0Ԝdh/��ȷ���v����Y���}W[�oA����K��C�9Q�x�o�j���,��]pC����!#^��6,��d���(���
��K�9�����T���؟��9��K������g�{���13�1��d�I.�i!Ay\Bή�y�����'s5ִTEEHL/��a��uF�D�Ids#ܩe�BO���5Q��	�b��Kp$�Ũw�[���un)^�v[v�74\m��{�$���wT*��#g�pW�����E��A	hN>��[�6z2���8��.�y(�I�r��C��R�F�"�$k0���dI9�X�:�n<=��|�n)�p��B��S��9�I��(㨙�e�jx�Z��O� SC�L}�}_6$���@�D�տ���{���N/ ��Z� ��q���6��5�rg�10�:�(ù2�;m)�"/xQeR�wW��=��������\�:���T��)�D�p�.YryZn&�DQ��,��n���1����50��č(�zq.鷷=q3�@@�"��1w_��V&�x�<��͂�%[:.��c?����s���Ƶ��{��{S��7���=߂�k;�o�2���F�N(��b!1.H�t�)��G��A�y!i�ODsЌX�Q9�\���Ri�:�3\���L�X��L�����xI^�U�:�+�P��Q&?�h������}��#%+�_�ҥ�ŖhY���� <�����b(�\4�!���$��G�Rھ4��(��S��rŖ�~��)��F`Yii�X���h
g�g��g|.Y��/f��s�_匡,�P�>	p�0*_�ᫌ�!�Sj֕�z�X�M@��2��O�Z��{��?�Qc|p�L78m��7��y��D���V��C9�]Hj'b8�i��|�8��cd��@�=~{(�Y}W��:K���
ł���]jH��/�ozQ�F�G��zR`엾�#����0����O�,�A��:�/��|��?^p`��I�4���Y%�cT�x0�v%b�}\�%�}�v�W���%����*4򻀨�m�[�o?z2���}�������?�do��E���]��� ��!Fo�r��2�Î�74��,~��!&��{�΀3�8��b�|�b���
>Y�Z�c�s�B������$�����x��mAw��t���W��O�L(ǹ� �!E}�a&�t����-eͽ3)�+�gj��v�h�O{�`tJ�;rn��`�U�sȁ��y-34����*+K˩t�[Ϝb�巣C0�j7�E1OB���v��3�z׀����Kz��պ>�8:��S[�۟Hdd}U������$�;Pe�%�=���N\�L�7Ep!�AW��f�1�h�%��])E�*��2�.W�rc�A�N�+O�����fE��s8�ao�ڌ_ M�;3�IIrq�[w����❱�j�����.��۔3�&��Hl�O.)=�|�Ø�����r�[����P�9�dשY�c�d�ˎ�a�{3�sG
�;s�����a,�b��������<����a�ϰ���(��J�kG�rt��Gŝ3X@.#f��%��FfU[w�s$,`�^7�?j2�s�}VV��K�*���,��$>��{�W��μ��\����RӢ��p�;��:�0ё~p�3U��9S�jg+�_5��6�t\|W�ڽ;W0A�4���X�NI>�φ�D� S�?7&b��rtL�>W�V^ �0FB��S����u�r��4{|��z*�^�y�&���mPrO��i�xBo�6E��z߫':���+8%���ċyj�_���&i����oNCW�rS̝L��DL�>�2���"����lTr��]�~��U<-�m���k��&�>�K�������6ȅ�'[X��|�!�%�C9�C�
U:\w�	;܊a�͍Qb����#�]!s5\��0lƾjN>��I����t�D�y���*���tB��ϗ�F���EC�#3M�Nm�	���m>�N���=b�]]�u��+s{��襕�:͂`7��pJ͚7�����sb����(i�E�gp��]�	��8��,�ء�zg�DmP�n�I��p��'��сT���a�<�d����=���"?�����Y���h�X�8���<RR>h����"�"i�k�މ��M��Wl�Pn�U��IC��G ��#��&�G�?����~��ɇ7U�Z�w�&c�0�j�����;��t���zYՌF�e���Z�?G���$:S��F�\cg	c+�^�L�Ql�u��/)w���Xs��0�u�g�`ů��b����^:�3��l�X����e@���k}޴�X�c�6���4(�%���3oc�V1�g�5m�e��]ƭbW�c�&������Z��=ޗ�v3%W_4�>+'���~��|��|1!�u=C*��4R���m�&���Èa��(��DÅ��"�Gw�VM�ɭ�L��U+c	S����o�����E�i��W2��ꝩ�� �|T5�_��(���q`�wIR;�kkg�+�b�lt�Ç6�1v�;j���TP@�?+ڿ{M�^��ٞq�B
��X$�WkA��-*��?8^vr1�&�&�N��d%p���׉!&�֠߰-�W�H.��0��_Fm#6��e�G9���8����X�7"6;|�S��~�b/�x+�m.�Cvt�wN�ɠ>��w�Uagg_K�FwӦ}-��`�l��o����<gaIm�k��׈:�o���'ջM�is�Jy��>����5�%�ʫC�SM����Aǆ{���L	6P�kW56�׵C��Ԗ,YA
�e�+�Z�{�%4�������2�)��j��<�gz�[�e�jY\Z�j�CV���8�ŗ��2/�6[�SnBW�:��0j�+.I�\)��άX�o��k�N0��L�'pRm�Ӟ>��9�z������n+[��i�ک�eX��9���+����1�9��z ��+>���Ƙ�nI���`[Nf�нg�E�����UUe�z}�����o��:	B2Al-���Rd�~Cr{(G1��ol"&��0�������˲����Ʀ|!6TUd����R��Gh������^��#pw�a��dk��[�a]:v ���h-��(�^Mk��-�J��-������[�W*���߀ ��d���1x������(V��Tf��}zy>�y���"*���z�4`ߛ��渵��^�n���E!& �gF$ֵce�3Cjg
�jl7�ǚ��n&d|:�vAL ]�U��<��L�r��ASL\9��v�hn>����j,
csL�K+�ׄ��\\��ފ�xWn��|���j�t���&v`��ﱮ��8i�!1��X3��/?�z[�����I썞�s؛�nv���궱\a';�**Y^�<)
|���̊5*�cW{�^W'�W��)7؀'��?h��&�D� q�_�I}���<�47.�0m��H��,���|���=� ����R#b����j��r.a!H�3������c Х7���J�9�k�#a����+��~�D���s��M���z(T��gXw='��������^g�{�Χ"���!�!���K�9�s��(��W�L��k,b�����{�H������0C'�xrZ�sK�]ۄ߾��YY�1�Mf13�=��ھj1�����p�d����̤? ��E��^�	�*����*#C�0c\v>�g�C\lJwQH�}��C�#�հ���
�	~�b����6R�V�����(�]�����0N��R���}�q3�kPX����#�փz����$����9�F:���p c�9�wS]�];>^c��x��)��Oo�W��t��2L]9�D��^���wl��U2��o�3�n
?7Rj�y��V�)�\o�E��8�/GȤJ\���
3����j���5���vPT�������$���j���a�����ی<UU�_$���}�W�����2$X�.���9���蔫�����/�n��1K�y�"����w�}�������,��+>l;�h�� ��h"|w����y��C�&���7��~�(�-�!���= _]قј[�W�̴G�bW�b�d\�y��ؔk^,�:�2[�ߪ�Ԥ��Ϯ�o�!�Rn�d{��jI�o���0ވ������,��j�1]_���A����"n*��;N&({�sw���w|��-�VJϩeN���;sZ�]�۹�o�2��v=���(��E?7�0��})F����`,��NM��"�4~��-]ʇM�EXK��V>$�����F:MF�����أ@�'�Љ��="r0�{j�x@��n�>'��/�c��7�_Is���g�+)]QR����ӳT����~����?�[���X�U������+�H��Cu|�m3������)F���0��B��1��?G4z7��tX쇐O.	�#'��ߴ�v!���w��i|&9���~����ː�;�2{2���$�J4:r�X�]�2P�w�<���=N��?淋(/<���պh�C�;t�˻M��֍o�1�sh�7����?=������~޷a��iC˃�����P�+�f�U$hˡo��u��k��l5vlQn�݄1�X�UG`v�{��t|�Y5��-_����2��r���}lDWr��J�{v�e���Gw��J�>������76�ӛ}:�Q�F;��ݥ�+i�U���3��+g�=���*�����6:r<>sʃ)z,M���_gs���������4�z�� J�m��t���7=���F����
�{��ë�U�Q}�ī.³A���y
5�&ֈ���;@ֿ��.�`l��ҵ�OHV_~�������V'��g���Уݒ	E��!�4��4z���|4��|e�>�l�[��:�G�����C
C�D��>j�[���g�`��qq������o�ew�>�yv+h�������ߟ�8g:��{</}A�[eN���6V4����a�;<���+��U����c�P�n�sbO�k(�E�o0�4�7�)��_��%���9o���>Nޠ)y����uzQQ�Nڒ��^k���vx�+�3�.e;:�gZ[9s}Yk�yq:��9'C�7���e�QWʀ:�N���y#��O�C���^+K������
���D8:��6w�
X���<�2p��;��_�D��,����J\�J��uۼ�WNN�(��E�+�
���\���2���]N��x=�-g��L(o��8H���-�i_�UƓUn�|�ɱ�q�*;r�l���A%���=SM_6�ʒ'S�9�Y2���N��a$�Y1m�gE�����[��Yp�M�q��uU8�:�!�����oԳ:�E��O��[���֟�oƔi8�5z����0Ą4TmW����grJ��.�d�����Ii�Ќ��	R`O�����h�a���6ϋy�ǂ��kt,�"t�/�m��1
�)�lO�uDea���u�e�|�҈Y]����wn&kgc�;R������T��3B+̾�r����2����w����[�]T6_4���,9����Wg��{��u�]x�H²���q�״.�M9�������v���O�n�ޫ35�L������uh9{e�:N�bE2��@��[�8S��U����Cq!���?�6��`q���9C%�_��'�y�~��QQW�&�(%ʿ~�Ϣ��=7�U���nb�e3IW�^��������Ώ��iM���k2����7���qڝ������gэ�۔��W9;`A�i�>/���C�d�]����'׋��]�FifΗM��]��%�_�'g���������To�@�.\e��1�p3�*�D���sku$L����*�֡v�S�_�-��r�'�.���I-=z���2�����M����T�]�-V�c�G���/�u���1�p��%��[!d�#~g������d^���y�[�$j��dEvď��{�e��yl��m+m+K�l>|��]����1���}�ꛥ��{���4����v>����3���H��� �7;?R��R�iߞ6�y�5�n`#O��(vc3����we4���>��w�M��9y_g/X����X�+g]Lj��J׹]��?\O�XZ�S��,��f�bg}�c�������I*���/o�ӿ�H�"�愺�+r�3��'οk���gi�C���C���{�������8%Z4��5FKcʫ�#	-4�ѯ:Z����0a_��}Z��r�%�.v�.9E#9-Ӄ�M[���u:�ʓ�R�`S���h�Ks���ƭr�r�����X?ֺ�X�!fT#�����H����������V�iץ�`����X�6�y��Q�UkПa�h�i��%�UJ�iċr�����ZC�nLA8���a2��@+�9��J�d�)H�ؔE2�tZ�;q�����^j��d&f�.п`�ȿrYy:�u�N����E�u�S�����J�]J����7u!��U'���.���RȮ����8)ℌc�ѱ�9�ql��Gw|�G�߯�����9>��?k��6	��8�yů����V�2,4��U����CH��!�7e�*�*wk��h���ڔ+b�0��w_��\F�J[]�0�&o�܂)v�������s���Y!����AfǕ�o�7�1o\�b���� +�M_P=��N��-��U��h������?��6�A�f�U�{B
	�HGN��0#1!V?��>_�nY�M"z�),e�W��j+R����(�5�Yn��AL}alFi�s�U���G��X&�;�����j�۔z���01p������E1W��ҝQ�
S���95�] �� �"g�I5��Kܰe-������k�����Z�d���R�c�q!� �E��O�)K#��0����x��Y�|>��5C0��]NDC�m@���<>�=�7m�&��b�v?�4�v.^���&(�Z��U"���HT���C:�GeZ�t�$� �U~��h�	��Y�`C�F
��ɿ9"�����|��ל���4a]��e�S_�&2?5B0>�d���pN������1b�~�ò_�_�Q3���I�>]�T�u)�?(aߗ>T�J����}jN|M\*�����X������HfPA�J}v�VO �������a��X҅0��h�j��q�Z�������ns�XY�eX�|���`M66��=�Β��rl�f㻖V��i�9ݛ����c�L-���\u�mH
�[�u"�ϜSZ�0����Z[ߨ��m,U�=��Nj�{�+�c*�u�2I�Cnh�>hl�Ǩ뢢�C~����, ��Z�9u�#��5�+o&���s���ZI7�S@�(@��T�5Z�a]t��À�V�T�s��#�U��zU���_D���{�l��h�|GŬ��r�{���<���f�H�"
*O#�?��Ȑ��F�����8�9l��^/,�h5 ��7<������*��^��i���#�VF��'���������f��OR�n�Z	b	�N@�ݠ�W��8!�.�� 7�=4eL*`���G�r`&Pn�4v@�	���`��Hjp�s�h]��R���bꅆ�&�KC��P����9Z�Z= !��/=�B̕�e@��N���o�V�%���V�w�_WB�CW�(��s-�wk�/,q�r,)�S���"_E�L| ��	��me���!M��mN'���ͫ7��*�Z"�L��������	cR�q���uI!�m"8�%U�!�Z/D_�����?��_�������<��/h}Y��Pt0ͤ��폌�]��]�J�	o@�5M�v�z2�y�t�8��Z�;�-��P�8�U{od\2`ΎH�Xc�ݡ� >
���Ս	��@�<�z��꒿D����w	ճ���4G�~�4���#��ha5zT��;wZ�ć\���MTn��m�9�r��Q�����D�D�j=Q����[cȇ������]q��{��R͸�{:���u�	�7�̵�����N^���r��� `+Ŷ���q��ﺋ.�<,BEr@g�3�)z#	_��7�O����k�E�ȣ���Fvv<�~�h��3�ـ�Q�rY�Y��?~\*O�IR�}�4� wR%_�gj��ߘ��0E�l4�����╎�F��V§�N�Q#�޼{��-��u���/�_HX�7!�e��FU�4�M�/���d�|�pl�?)�^�ҧ�Q.�n)��_e�a[�n�v��y�$�^�/�eY��I��@�S!�H�E�%�b��o_��H>�*�3�E�Tg�;����T(5�~���.�"ka����_��kze���"�^�Z_"DL�/.y�ov@��Li�p�|��}8
�Gm\�ř��2�{hFi����4��EA6�D�#�|#�ۂ\[Z4���nV�h�~`T��h���;$�̎�+��F�í�e�c[��1��O�G�.A�.e�x���k������K~���n�Ʈ.�4�������'6/��6ۉ~P}ҝ��n��" K�k���S�j��:S�?����h�X���M��?m� {t�MR.�_���	��VF<�??n�\���	�����S����Za�H��ȥz����pj�I���I��|~�ٴ(JU�ȧ��,p%�Ȫ�f����l>�.��A�OH���
�'��6�ȟ!XI}�}D[&�!�G��v�ѕJ,>)�^CdG����"�Z�E�����%�`��R�[���doao�l�#I�=p�qv�YI��7�U��+��t�ѧ��&k�c�2�BfS���uд��/�A%X�� "��ib�ԣ�߰�uV���e�	��g5��N��������ev�*��-5�=%��5��\�-� �{��hk�Q?_��{���f��d[�Qta���?�hjV��a����줌p8�� ���B�_]�K�y\vt�O<˅+��&\I��G>gH��-L�K��/�[���~�h���	����y�q����铙S�y�wD3�eR�48��&.Ub�Q���>La/W�%�ڙ��k�Ex:Hr敗�{�{bѻ�s��]"�3c�]"��q����=�ԹIv���d���=-�=� ��b�~��Z_���j���?�ld��+�L|�ѵ\�k� };�o`���ƒK�6i
i�p������Z�J��*uE���s�y�K���i��c>���+{�}�}���O��W�K����y't/3����[�r[��YDeU�R�r�@%������T��/���c���l����f���e���BqF�><B���%��X[/T"�G�@�5P d-5�5d�e����w`�S��I�G4"���4Z/?�j��Ht��R���yF<JV̥���f@�%W{�w���=���;7�8jG^�v�
Ww�kv�nH�|���(��6!���̎����pn�� a��f��(��?�
BE��Y��&���'�0�,��3"�jl��)�o��E�]��'!:A�՘�R�*���D��r���p%5Q���'���ި|m�L�Aa�7�ɘ���e�e��_@�&��9��}ܥ����=�E72���;ʪVB^Y��4�q�v\y\�?_�&@�^��[��۳�Oyyo=x����^(���WdeMBBBN�w���ݽ��,,�**��u@\\|�u����ٳ�o�to�x\VV�6#���d�葠��~RRbo/I�699��B2;;{/�$LPɈ�,��|��i� �/#]����NY�qw2�1v����|�|s���Y�5�U׵�Rqr玅ؽ؊�[6���U�=��L�ww���s��q4&�H�sg��t1[�=������r����t31�gO��DS���)A~������Ү�oLz[!nӞkQ둯����K�?�I/jm5��?TfcX�dY_����|�:vv��!�W�.�%�X`D�r>}�"'g�s7M��c������,A����4�hԄ�v������pJ{��d�L��+���+]�k׻>�Y҅Ui(|\z��8��¡"+�J�Ʌ�b����z�z|��d�v&!���U���эH��M���h�Õ������*u�0Z�5~$��C��?L���&ߨ(��q�a���9�I��@���2Ft!C���w���1i���Lu���ٟ>%�����:�fCg*�lGK�#zy�b��e����R�o��љs����p�Fi �c�l>Z�R$�۞����Oj���`���6{�dl��t��;L}�oI.a�	�� L�Wzy��/�ut)��	Ч==g�Z��2��rdDv�0e���Ea�6_-�=22R���m�1�xWP����Qk�;s&((� O��[C;Ez����3��f����.E?�&#=�8F��'O�p���{��#������ؽ�GO:)ܱ?���@ļR��{ÚX��2��BU�޶۔i��N���
�J^A����}�v���"��eYw�d� oV]�@ ��(�卥��2]��,,.�^��Ū{tvǻZ�_މ����<W���+p�.�����Bźi���r(�� ��?�?f��s�G���,|{}	�	����UR]�dݮ��rW�����ڕ��-֑3'���Y�锭Z���ҹ�E?��Ou윖c?���D⇌��b�τR���g��u�# /Z8���y��ED'�x�Sm��LC�$e� ����E&�����o'Jߑl]��4M��&�����o�U��C����P+ۃ%d e��+�GA�EFF���̳\\��HģG�����с�U�ß���������O�L�}K7RG3�_{G�?�}��������]�7̀�0���"D�R�͟:��'�l���2=f����c�����B�3�7����w!M@ڙ��z���Cٿ�-���
%��RYr�3�W2�,�7d��N������G$o�Ĝw�g����.��>Ԟ���y��;�|�@"٥J�����y�{C�m�7��O@��J"�K�U�c��������:�`���.��T
]ZkI�Z�gYG�w�x������AF���8Pe0H�(M���ȟ�)�cw�lEL�w�6��-�~�ps=Te7��h=�tX�{�O�MҥΖ7��N��F�,|��`)[]�<�=�b.	� �]9��Jǈlo�;��ND]�oo��x�J���h���>�3H���[�S�A����Fqy(nص�pn҅�ߛ#�� +�������6>%O5�d�_��������6ݗj �3u�}�c�2��S3�9��_|g��+7f���0�����|S��Ԩ�9��<�	\���Tak��,7��]��fƎE���zB��2s���k���^�9�ȭI)�z������`�#�--��Ė�/�ݾ��d����{?�Ҏ�Z���<Xrc��u��v���FJ�1����������6��;?­�
f��6e抄h�sg�N�Kp��%�}O�I���˪�V~�%����wo�3�/��=�d�F�Zl��lQ��|L���ո�@3QЋu�K�O���52k�z:�6C�4���Zv ���U)�}�_v<vJ�#Y
Wf���^�کӧ+���]1��u(��S��YY�����)�ii�kOa�C� <��)��pծ[8	[���ev|� ���	�m�n�<V}5jZ�b�Oѐ�\�.�����f���	ƛ0I�D��1�{��͌�kg�oצ�/S�rcN[|�n��r�м�xET"�7-y`���O*�M_ ��|_�t���S-��G�����<�5�<��$>~*�+�?<�녘�_m��o(d���Dz=N�~�HT����1��/��VE�
�ҕ<P[!�@w��|"��Fs��v����� ��OCj� ǯb��&��a3O��R�Tǥו�.c������.�&6
�5����b/��8!c�����?U�Qt0��
�h�q�7p״��qq!�mm���1l�I��x��f�pl���L����[�3���[�o[��n��`�O�T���zb�EPӕ.3 ��� JT��ׁc�~CB�7���:M9x�jCe��h%��i\���r콪�#�$����z����Cw���A��a���l+���kA�Y"��0��]�[�-�w�p4u�>���U�3��Bg��k�O]:�P��!����չ���P��הm[�p4~��cסsK�y�n�L֙��Q��c��t43p��R?��Y�7�r��y;�t�^�F����k%���d�����t'��Uj#�<<�D�0����ele��A�^y�no,G�GE�ߙ5�.��}��.Q��1�5d u�$�;?1�%�U_L����]��TO�o��d��h��'\x0L��q���=�̕NZ&��'~���;3��kW:p5��։H[jjQ�kU��@�o�s�N�E�[Z��K�-�w�ȥ�j{k8	�*�;&(-m�4\m�"�����@��h}�ر\�LB]%��˗5��qԱPdsӰ"L�9�f���:{��5�a�z�&��%%�����/	���
��w�<�rT�(�c��s<{��rz�;ub-Ce t�V��ۢ@ɼf<�\����g��a���g�1B�:hP(a]�Q�:ZE/�5�/��l<��PPr��T��'�>�N1�3�}�V
]���9zԻCj`�M �/U�S�c�7i$i��/jv֎�4l�ڰ���λ�55��Ef8R)�QB�%��!ʝ�;%Н�فQ�v�z�m�%ݱ�u���&�'��,��hT�dQ8�����j������Re����K�O�O�h���8�T�5V������]�h6DZ(�Z�_v�B�KVPt3;�"�/Amf�Yk�0RS���+ߴ�v./']/����x�F�<cd�O"��o�j��ˋ��̈�/.r�Ü�\���SYl�'>�,�:������D�B_�Q;E�܊��K��*ޘR+`
�*�93�d�ǹ�+6�qd[�p�����8�x��f~!�J�@ݫ����5��U�
�35w[f�Ք���o�����Z��m��D�rvJ��E0��,�ޅ~?��֘�d��:�X�bKp�� �Z}E��7���F�
 ���l��y��h��Ɖ��K�.ev<M8��ؾN}�<  �]�ɮRE��R��e�3�����d?q���Ý������[d��U}6=fҟ�w�x�Ť�NW����tf<�a��y �����Yf9�*����Ӿ)>��^����ܹO`��߉%�{�oo,��+��}����Ѓ�G٢ܶ��Ǉ��wx�k�qX��E�]� �[ì
}���β�-�u\ɏ�=�н6���W'�J�:�,
�a�q3�3������/�gO����+H�ޑ�b�G��O������s�;��z�]j�|b�T�8�Le��Hb"��*L�c�n�5����,��[�֫*���C�q��`0fv:�
,Q>�f���D&�ty��W	WM?�S1�비L��lH0Isg�6���	�ev�S����k���?��9���j)�Wb
%��)�EIK�D����s�$����i��#c������8�+k~N��EШ6�4�aB����w�PR�]j��4~������.�!����(�̥����ͯ��� A/��|O���=`�Y��]��a���vk��͉�v-���쭿Y]��f��mF%����o��^&V�{G��w]�g�6�Zಢzoz"�֗l���+.�cB��G��[����݄�hG��:t�=o��M6�W/���56��p��F�jJ[��i�j�����Z�����^��m�B'�-PG�A�n��n���@�8M�;�9HG�V�% �Ǌ�?�`�J-*	�G���~;"��>b"ԧ�gB��p}�7��9�K�����uk������ Cc#��^
�:Ke���,Я(Dq9 ����Y&X�Ch�֭�׾��B��+CJ��g/^�t��5'])�a	_��X�U貖0R�{،V�f���!����xt�;�P�:l�K�TP�cN�_����,�x��)���}];����+��1����z6�Vzw�֠s3h��x�O,�ex�oo�nX�'�i�^���0Y@�|������_d��������Lu&ZZ�!�s0��C�~ ͔ev�ۛ����\!�F����,£�c����Kѕ==Q��OKi@�^���~#�(a���Ӡ^{�T$��)�|�HA�t|C�'��Fo�<=���f?���vE��[ P�W9r���Y�����v�ߓ�6r��\�>	��~��K�K�%���Ɯ���x��GEҜy5)E���~�9	-�����qǿcه��ע�x m��Uӕsu�W�.+�ݝCG�����B��;"���B�ߺ�t�JF&I 6�' �J�D�m�M��R�e�O�C��;w���U���H���;�Wܾ�WȀ��(��.;	��!�����D�k�׶�ї]�%�~'�Y�?�},p4U�O��\����/v��f���0�	��-���=�� �#"�������K��߾����*$&vH5��+�<�I4�t�6��W��D��gңb�Ha��� R[��+���M�赹�ܜ+O��cۻz�̕���# �/�O��;�a�-$%�����y�!�����'�����M�M%���;C	�� �M{�ƷF\��w��ɵ�����?�ό�ASM	yzّ$Y��1��������ecբ��'��NV�/+F��6�3�`���#[:U��~�#�)l��ę�K~���_��/�K�>�48���~F*���C:\�[��/�&Z�C��l�OHD�E�=uAn��0Uf15z.��ޔ�5eM��
^/(��z��Gێ���VIg��7yԒ���'���žBS����)�y�JnG��� ��z�>�7��T\���m]-p����z�\�n�migf�0)�F�>�6*_�_�9sCj�4��7�~k������O����>u}�]>�E���J��:Z�A���n�n��2�����^C��˽EWޗt��:d��_p�v�^]yFF�[Ӈ��X:����Uju�x�y^������z!�L;!P}�@]�0�7q�y��n����*m3���s�ᕮ?��?5peX@
 �'��vp�:�稖�7�@k&��l��A�q54�o� ��`i�J�!9��D�76��mR�=U�e����Һ�bT_�3J����_���1�:�������e!!,Z㾵���h�����I?�oxV��ߑ�I�=���/�zk�Wl%�ү��^`a �*�]w~a��S�?t�]:�Va�J�ߪ�gA���~Sw��%���}@�2�ruɺPχ��7�N�����O,d�Du�VJ�]�d���ۡ,U�Ǫ�do$�z�Wõ(;�d�[
	�#���-�vu��|�p��Z?; �������h�-,i�>�lew��cP�R��c������d��4��l�[�8��b��o_yz;{�Y���z��ظ!�|z��&s��ϙx�W���^��911;Pa��W�h���!lc��#��|);�6H�� M��֗/��s�_8�u
a����f�1�؈�s���U�Xt��-�ұ0���\��d,�f(}I#	��[�5L�?U����J�쌐�AS�TY�D�Oa�.��ig�t�IĒ^�s~����*t��x����b�9z�x�y��h0����9y��|f���$��wI�䨍�C]����-C[Cf�v٥ܚ�w���yU�7q!�FLak�iO(�%�~I*/�,ZX��2���M��tXmosX8��6�1�9 �77��@At�5'�rK]����Oa���C�-�R����덙�˂*?\I�?��~�$@�i�FXz�qW̱vk��R��=��{4�.��'���_�|���Ew�&�<�x��0�ܔ�$iCa�n_�����@�fW����)e����;R(ߌc�J����? �		���!��� ���]�)7�:�T�~��NeA��:=�x�|��7r�=|�=�=Z"^�p���*N)C?��8I犓��EÆE��x���n�C��7�8� ��H�:�Ku4n��z�9��VݡZ���8��8�O���Z�p�9�q��&�!����o�Z�x���B�̳���Ro�o;9�k'gE���L�Ǘr²������ ��ir�RQA&҈]"�K)+ko�ٮ�rU$��7�Ep	�#�gjB�n�����g��u��2���]�2��ng ��"�ݰ��X�,�)�0��	��J�V9�y�H�^M��*�U%�s� ��0��{ ������q��xSPP�1Z&�f�������+��]  �b,���l~V_��vWW� ���)�(�f[r�,����g`]�(��s��zvR�dF�C�U����n��_p����������;�b�xL����C����XD���o(��ӣ� �R��@A��S�)Y�i�x�^��K蔗 �����@^H@E=�����"�Qf�C64
I ���|Q ��� �B�x��)���`\)\];C�X��@^XvcEB��G7	�9���{`�ۢ�;�D��8��^�P� ���'�wQ*1�q��?E��p���o����.���bCA��S���Uo�U���]�ZՑ�����(u�Ń����8e��Oh��z�rhm`��Sy�3���o�&��$r�I}��q}ĳ˞2�K�vN��QqeV?��A��\8��{	�=����>`7�8;qdv8������4�{z�wC)�b��H���g?j���y���K��RH)�b������/v���5��Ƅ#d�"& AW�w�؄��;s+���F@,��Fj�A���.�4o-�Iy�Pt���.5j�!��;U�R��!ͭF[�����: �穇s;X��v���)�l��_��:���������b�q'��Û=���0�2��K��l�����@ �g����=Rc X��ܰ#���1�z �[�Ǐ�W#?�I�hT$�{,L���
�8[�q����w�b��Y���w�<�zW؈�����k]~�v�85�y/1��@���;����{-g^����p����.,G���=hL�¨�b�@{Y6�3;"��D��~ �WH%y��`�`;Ef�]�;�@ge��oW��C�kJQz
�a��\;c�A�?1A@T!�����B�����Ls�g���(d��£~��J���M��k���GT���_�t��G�fȾ�C�8k��v�������r	DX#٬ڥ�+U�. $`QЬ7����fS��
����h�s�4XW@]soKJfb4t2�"�xƜψ0�-����#+�`����)d��f�t�]�\rCgݛ�K�.Ł�6��sSka��˃�W:+1�X._��N���N����(���۳5�QHY��w���!%z幁��͐���΅t]��E����8[�z?�:J��5�:{��	(|/�3����6&`3Ф
��#N7&]\_p~�����ɾcB*�"�B9��Y�_d����{A)���w"����
��&�r5���B���(pYXc���o�	d+eGt����E-]��}��O����]cL�Ւ��@*�mx6GKK��K����4���ƀ���[l�/�N[#��}��]CG^�UV�/�{�o��@��4yHA���������dY����0�Û�%(�����-P��􁁆�Yb��J�S���ln.�Z
���d{����o1�������oEbM7?��l �c�_���f���;N�ǔK~Ҡ�j��(5|(U*D�����y��*�㮼%�"wv�0��G�@��X4
\dr�3i���BU߀ߋ7�9�����2��J�Hi��#�Y��@X��	X���]�j�A�lW�tk5t�me���foYo}.Jڈ����_�����f��j��D/��*� ;��������(�	�Z%.��U����Z�kǼ�>d��-3x���/�&�@S~�;n�L�F�Uء�`ˬ�%n���AȦJp�v[�mL��/��ɾ�����?N�c�a~�R�����0����;T�.������ed��߲x��pI������$v�a[�d �r�Ĺ��:lG����еQ�2gg8�H�0�zz%���),u���'(�V�h�z���#��"����-����� 2��ꬪ��hL���.߱��(��|�<�S$G+zL��<�F���T*��[��R`�gH��sT��A���" �3ѕ�g+hv=D�v�͖yY4Z��;���jM���6�۹�o�i�"2� Ѝϰ���%C砵����ԛ?;uv�GK:�L�3�7�.��tD��I�`~��x��� m	�Zu�|�i
�y�)3����	�֝�)�Z�m�@��a.����p��A8~�<	�Q�F@����O�U��1�ӑ7/r�r�
�ޛ��ݮ��63U�=�Y�?\�,��Hʾ�XE�.쮴R᱗����5���Cb���m�Z�e�mu��C�G��F+��MV�o�M���y�k��N�~���v˛U�9�
9���4TV��x�_��#CИ)�"�W^�ߐ�+]7=�^��K������d2r��ҹ���aaK�BB|����6N@ϓM�3EK3��l-@���`ݿ���9�Vݓ,����v˄4Z6糇�uv�o�%FKO�A�w��D3��l�s����&W*���[�ߴg�}ˮ������_�ըpKU��Q4�B$Z� ie	o�1��V�9�fu� ��4?�wnW������߇�B���gvL>�6��
u�hH4�&=f���1C�	�ݑ�>��je�	X>P|�ek�8O+�y�{�,f<��o�K?Q�o�nAҾ�����0�'N�xu�fM3mؚYz���]'�~�e�J$���N���l<p2F\f6��H|l>tu��rz�0��ԏv����m�Fj�AT�d��t�v�ĭ��V3�����C@���}[�1�q���~r.G���W��$���ɓ'@ �8���U��EAg����M3��Z�Q��}*hx �R��7wz��G\�$�ݚA�etü70++<����=��86���YB7�b q׈/���e��0=�C�'��|�f�������gB�d���R� ^����Wf��� ��ʭۻ$ĕ�?ZM��=w0F������ݹ�_yb�1$�j(j�Q���e�	z3u���N�8p����;(�A8(��S_�9#_����Ά�4�w��O�����(9>)�@&P�[�Z�}�Z�z�.�p���]1��Aw���=�v����s'�P�]�_W��}�~L&�+���>BO	|k.f����u�/���|�+��Wp1��p�mG�]�7�18��^ �Ik�����\������ �b�<.?ݥ����G��a��KÎ�����e�L�۫�����{Eކ��(�]k]a�a��?C]qr��15;��j)r�r��NQ�����2���	��,>Тo�l�cT:�o�d�]�3���
r��/]�Ce�}�P�hy���g�l1t�J=� ���770l�Ԍ��FDW���-�Bi+�>�g	�X�fG�����[�lj�N%�Z3.Sґ�o�� �HpLE�:��/��~e�kK��"��닰̎�T�J��Ol��Ŝc�g�T��y���В��M�T�F��甆�L+_8xv�y^[z����"ػ�{�wy��U�\B:���ߤ�m��W�~�h��Ȟ��\b�r�m;s�Z^vS:�]����={	(���G|��Ĩy���8	Å5{
V�n,"�Kz��_uO?=�,�&�|J�t4��4ˤ�zY7�ݺ 87 %�6��ɿ�oG���e8���:i���%���Tk�Q�qR1��x�� �ѕ�w�X���P����I��N1�����>���(�w_���:!�9،8r�H��|�s0�}�!�q����?��v����#�z�g�3�hi�V^yr�5߻�9/�׫���,�4+xx�:����[�_)<}��G���;�H�ǏʨAS3�s��{�gm]mUvv���u!�I�H�hZ齅$rhGG��I%f�U�!�;�X)Egt�-?]�A��ia�1�I�xcsV�E��3�s3��D��%[�c��E^��w1�
�1h�����NU��EL�z��z�\� ��n�ݙ.`6*s,%��#X���h���o���{�`��ƣLZ�f��5�x����s���(Zel�⫉p���K۝O���|��~���DZsA�����4�3ݗ�C�O� �[�7�*�9�`����~4�9��C���]=�T�2m/�]}������)��_lR~�u+���P����A}p��u�4��>���w��K����/��4g`�\�#b�+����$	wiN�y`�zNrP��U,�?�"�_t7��lL���)�W�#u�L�;�����Z���G(q�kL�i��9��ύ+\���]�w��wB�#FCw
,:	:�4�b%>(��CJiJr�d��蝊�-��pϭ�D�h��>��{/s�����ʁ=��y��eM�m禒��I���O�l	��ݽήoů���9�����8��9�L�E��]�~�7U�ؓ��M���l5�[A�?t�<j�9��u�1-d�(�}ĥ�uf�0/�^tlojw+:��M9+-����
=�q:m�zL�����g���6C]]�S�`7իG#[?��<���R�Æ�IF��W
i!to�KFS�f
Aj�pe�Sѡ�`��ج�o����&���Ɣ;�O�8O3�o!�6�s�T�N���X�B��0���"�-|{��e��qۭc������������,�1?��p��>C|�i[{�	�ߎ�x_�׼���%ճS�����;���)�l搮�=��c��]������v�)�=��� {"��~�1q����G�K��~��͟tO�H�_[z���qCol��R/Y�2��cu��~*��J==0k���v�0�ŝg��U�X�.��u
��6� b
���������ʹڭ�-����d���l�����{[��P�Db�YB�K}~>B�?��nG�h�����d�l�a[c��~Z��2�S��mf�;��r�U)���m�]J�D�[P�:2o����˒��f3c;锗i�5/��x)�9���3O|{���
��u�}Ax5�9 �^������ �)�*��[� ���WWv���j��<�,v�8�)i)�(����f�n�Kt5�Wo�~|�|��\�o�2]��B.�P�?��Mf���ΆH}���'O�Q�AM�!�y���A�{���:�:2?)]_��l��u`R��#@>�c�a�e�H%S?'
Vh�v���V���b�����|D��ŉ�U��y��V������B?-/^71�/���~�d(W0��;�J���7�#l�s/*@���c��D+��4��w�O%Z�c�q�+.,���>��`׌�ݵ^�N����>�s:�MCzC~�V[�r�@FhH�]�@���F���$��I�ʦ	TuP�KϞ�@�o�:&�a�M�C�Ii�*���Z�\g�@�@Qg�lu>�E!h8?R�־����:�t\^�s,�����૥��W�]"iGN?櫾zy{3��ҫʓ�����+4~C����z�ԯ#�3ӆp+C��a���������q>f0�ˋJ����PR�H�����nZ�6��K>pI����ur���;  ���q�˵ٚnT3�KK �ިl������:��ٝ~���"�����w��5RQڦ���Q: 5��麿�X���O.P{D(�jMV>�x��6��D���2�\z�-5IC�mL���F��	�E��|�6��\���VԬC�k���v�,��P�u*9�P���b�;�沇�[�@�uU�����G���'��d5��|�QџtW	^���4`���瀞����1�ς�@��h���1%�����`�[��ǘՐr�,L�� �I^��!�R[=���#�����Z��z*�?g����b�["�����=��sGM�1U��b�a���f���!"ɡ��Wp;�#e��|�s�)�Ц�.�sQ��
���wS��N�Y�L��v ���Hx&=��ǯ���ٞa��U�C��Z�WJ����ø�~}������w�.W~hī�E��dnמ.Ҽ"��f�yP�o=�|�����~�Τ~�|���o���Ni{o���� ,�GZg�����%\H�	��u:J�-��D\'�ͤj
�T>�,4A_�m'�.��<֚ef�0�q毎�;/�b!�^﹓,��V���?Ae���Y�y��`�ڜ_�W��<���ŭ�(v��:X�Iyg����So��4���k�VU�:� n2�E���@���R���6����r������t)�(G̧|_�����7����'��R?�p&8��dI:���z�X�2Վ���l�=�l�]�!�2�����i�s�:�������!��'%��j�����7��0�����J�z�����/=�a�kf�}}ɚ�g�7o�5�*���)�f�ͅ�B[��?�錄a�(�L���θ@�$$T�	��-���c�c%yx��̜lt�Ue��;����䋙��9�d��!8JI����E��6)�f�ĭ����ӗ��]mw���)������(v�+P_�L�7�8ʫB�E�T��]���0�|�0DڐFȻɡ�?�3��1����������S��ٖ����� ��!��]���}��	������`vW���k˰�>?���D�WGE���yk5c!O�[�@B������%|������@a5Zk��u���_bM�G�%��6Y����(����� %�`{��
^Y�Qj)2H~R�M�flSN��Vq3Ri�D���!���,�/�O-��_f89�qIb�㻺��>�_�԰�$$�\��N7�9������n/X>�$�Nz*V3R��^��J|��^n��ǰӠ:<�����9P.�/b�kuP�ض���u�Ĺ6�G�Q��A[톪��nF�j!��<g�S;kX;Q%�5h�Bs�z?3[�����5�7�׏�]���ٗ�Ӡ�5 $;��<�3�ݠ�������j!�ᢝ�o���h�o�n{�0�.ή\L��w���U_����/�V�ȃ�uܗ�)�媶sgT`젙�ظE_�kZ各�q�"��s2$g�g�@�5Ջ��v��$"��4"30M��F� ���8%�Krʻh&��Ar�6y�� �����M���Չpey�J�����+������#��Lj��nTUC����H���R�.W��j�d�2 Kj��Æ��Ĭu/���/���b���I�����v�a֚z�$�e=@��+�J�qi@������u,�؀ ��|-������ʖ�4����nB���v�X�H�ƛ�ױA�h4��\	�T�?G����R�ڊ���+�0Ih����Y�l����ء�a��./�Ȑ�8(�3�$��ԥ�'ng�3oᎹ"����c%��1�W_K��Od�����PZwİ��P���W���^GXpC�I��W��=ݧ��[c��-���-o�Ҽ����濖2"�������mjEGJu6U������W�W�F�Bt:
�o���+C
�n��&�24�p+�_�ȥ9ꛏ��x�z����U}���Yu�2J���F9&�g.�SY�!�x�cQ���[��w���)H2o�۝၅��-UO�aE�����͏��'_����u\�RM3�M���ϖ�� ]:x��� ��3�3bJ,�������\��ԁ����nO�}Ƴj��(\��8v�8�`�	o&�?��`�lϙ�-\�c���~�i="��q#�/�����]�&�FE����FSW�;\�S{{wЩ�a�	׹��:f�t3Swuu���s�&������k�!Ҽ��7ǁ�>4�����?����l���`��V���D��uE@�"�A�tU�QAC�"E���
H�I(��Z �9O�����g�Y.��9g�����\(����$��Ӥ�3�c�F"��K&^����!W��p�,Gq�#mS3�1�XVч��N����C�ǱsڒO3��f5�d��*�*=G�V>qxd8��(_�J�o�����!��e��]0&�/��}j܅B�����,0`���"A�j45y%�W�����<��J���#��i��N����,i��|L2Ɏ�/��9���%�~�{G%沦^ �~#�(5��q`!��<"�u��V����h:�������)���fQ��"i{����\���v��0��?$\���$H�,B���m�ʵ.�p/.�kgkp�w^��~T����#���%��vǾ�Tz�l~R庅���GBW7l̎{�vw�Z#l����2��r� x��y��q�l9����U�A�#�5S��W_��η%��������C���2ݼ�V�4�ۡ�j�%-q��0���`7Zr�ښVSF?~k;�>�);>92��#�(T�S���^*>�!����3�5��j���*�"��%R��(���&f7�Aq�%�Φd5V��2��)�U�$�4�i��/F�s�@64\g�n �,�X�:�tZB����|l����L:�Z(�;�RbT��F�uT�/�U����卣Rǌ�H�w�8G�̫�ٞ)�,���e��� jv�~jsD���i3��M؇�H��r�l�3����j��f�ި���򁪥}��a�[��'^��N��˹�L�����:O�Qe�^9ְ�a�`d�dP]2����k�;���Ϭ��G@ݷ��l���ö���GQ���0���0����w�����\(i�{��X�V����$���	q�J-���l��Ĕ�n�?7.���w;��Z���3���Mn���i g>��j��z\��M�� r�D��/��ޞ��ϱ뵶�DE�ffz{zWz��+��K8�d�D��ܧ��|qZ7a#���]ZZB�ʅlI�⅃�.3�dX{k���~����ǯ۷O1940>�^���oFz�;r�6^��N��	ƩbA�p����Juɔқ�`���ڵ�i���	#�6CZ|a�ъG ��&�����v=g��$F�r�d�U�j�P"Q�+SS�O��}׎�{mϯ|f����z�����.Le�Z�\��Unp!|g47l3b���d9@�|Dm>
[��ZcBV��?�L�0U�ha��]�`�c�5�2��_�c��cq��W���Ih�J�N�0�È���UI�\��+�m)�Β�,�
MW ̐X��J��$��c��
e��f���V�iE��^����^#U�L�����#�u������C[N;|)S|.�I�f��.C�Sq�^��J�#;	e�Z�^ t�K�'�p�����;������E��b;l���5nV9,�V��,�[&����=֖�I/��m�qzU[���D�|!�Uu̱�oI�-�M���pc��.?+�FGHq<$?�B��Y]X�#�KW,�_��^�|ofX�aǯgj��R�T%)�cE{�q�)]]�!P���|����X8�����+Y����0P}���vi�[�U�� �:�w���a!Gj�`�/&�+,�0C\j��y\�?^d�E* o�zO
�Ia�ö�ΡZO�(7a���7t���a.WQ�1���)���O(�;��Z4��Y8J���{����m�gIr{,=#M��ujJ�W�Gv9�2]�*fr�
?F�X�dˑ{��� ���*�a����T��=z��#<��[��$����S��'���g�H����tT%;�������SJ�=��*��l�g�����\������n��*��Kr��^���.��r�%�К�  �t��@�m��:���E�P/y�0qdg�b��Ϻ4sy{�)��m٘8٭P�O�i���>V2�X���$�������O�k�`�&���FB��>}�{����֓k!x�hD�mPW���n�kB���.
E�0����w��Zl�q0_V��* �^;�U��1�"�nľY�����g2�����&�>�)�����V��.���s���Z�JS�?�+5a�"`�zsFƨ	��K1���q!2��ql��~�������]��v�o�nb�^�uI��ʁ����X��'R?b>�a��8��&������lg�3??��FT��A�/`>�_�� 7�D��^]�(_��a�P;�A�*�Ja\�uQ��Sq�����|5�je�7�@��4)��狿u���U��F�����-s��TF�Ď��j��x]d��m���m��zc�z��ө{!�q��px5Rܬe�����)���J�P9��z�Aٮ�U�˧KV��jM\p�Z���8�^�+`����3���^��<�-�k�o+.(J�7����(�������RC�|��\�]G7�[��˚�Q�ӄ6&P�Ck?V�ksfXB JSP�?d�ݢ�m��k�
N�n��{5����h����$�JK7��d���h�fT8GK��X��xj�l�{'	�6���f���m㯄�Ш֟���	��c�u>}�ϼp���9�՚ 	�zx�n�uE�Kl����LHG�UB�AC�|�K�JL�0�F��z��Jl~��3ʇ˜QA87 񲜢�4H�ꝓ���1�3uG������R�^!���YE!q.���<7fq�hw�|T��[. ;$��.�T��2���*����+��2�nz�u�B��Q��#zk����M�ǃC��f��a{���n]�wv��v�����5K�i��
�:� ���9��g�5��r�~�����i�\m폼o(��2������a�����<1�)o��H�Sr���f�?���86:�C�#B|�M��s=OJ�]P���R��R%�O(U�o|s�.Ev.��t�X��J�ſ���/�߇5D��{ nA���$�B,��E*�307��@�r�\�?����*��7w�ݏ8�JKK�q�T�)�M\���dc;[�h'�su&�Wjm"�sEY��k�t���6���[p�e������eAA�*�N"
u��J(� ����Ж�o��/��� �y��3�v<H�-(������9�P�$���0ֵ:�@I����GN	���$yc��L�Bq���?���2nj���>�ŀ��b�>!Sf���v���ԖK��/oSTUQ��6�H,_�XP*O�'XMV��Pj��G��b�� _�c�
���B�<bg,Ǳ���{ۑ_��<Z<(��@�������G/�-��(C���X�.�/[E.�q�cȱ������]7C�!?1�O�Pl(����t��v��o/��(Tu+0���̯|�^?(�|�-����COr�塈�FRJ�aws*%�F*%�r��)\5#?T�|{`0!��'��p��a�>6�,ws�P|}�J@7��m�:u��HKPf� ]� ��NK	��T���~N$��S����4�\��
�V'_�z� A�����B���Y�C���P�`F�����n����+���s�{�b�Yf]_^���1Bء�B(���)}5m��fST]�,v��C?�
c��S��Mn�z�����-�I0�
/�z-{�%�u�3���[ˁ����oH�P��M1R�GO�_�����<p[/�)�EӠZ�E�2�Z�"���]�J�#EC@�[(�����pZ���"qt��3���h��J���4t�˫sc�w����q��y�i�Pm���79q[)�j},E���Sѯ���*��5T%.s�]B�nal^榉mT�w�~����\.\_H}���Q���"�)'z��B�Zd�������2�* �Nv����76UK�RͽX?��1��6Phu�Je�:_3	��Z���6�[���G�5д�nU��7�����]��0uG�~=tÝ� �K��1%%�<��W[Zn?�uyn��;�{�|p9_}b�=@�@6k��}����g�E�� R��*^S��	��fwD����A�`V,�O<��;99M�嵨&���@�\�cw5&c�0+�o���C��t��@�&������:���Q�ݦU=P��{;V�J�@�EZ�ƿD�2� ��@ 9D�� Ľ�h:z�-Ox��<ƹs�e���L�	�װ�G� 1�yXiɧ��r^ íHLL��, ���Wt�e������*6����ٳ@���+�x؊�aI�ic�I'b˯�D�#7��>Z��O @�`x0��y�ȣ�H4$�5}f?��A�;0�i[_m-�,8�erV��뀝;)XG���g��c����k5�ss�L��;�[:,�o��G���zN�;z4����D���̡�٘"Q1��`O�|P؍�-0�0��s}}���W���U��|�L{�̍��}��ۓ�)w{9��v�s �G�u��,�c��%�2�P�oT�vV�g3u��U@�E����ُ���z����h0��r0���	K�30�0�j��3��M_�E�)��Qc��*[ �ص�,�ޚ���v��	L��7ܓ-�X)�*c%����)�k����C�؁H�qի�Fv.y��v�GX�a�W��a�'��s����?�������Y2��r/�7�
%?F~�V�T`8'��#E�E
����u�htiY�Jp���j��L�%��D�4#�޷���5��V�c2��/9��^Y(��pv/V	BzEJ\���YYAt�2��|`]O���b5�I�����pV�׾R��԰n,�a\�7hc�����9[�+���Q�����Aڜ+����(��������:YH4�9Jfp���ʙbyQB��k�I���8B�@�"���pN��`x�%���y[o�RI �a<ߞ/B,eҘqą�I����-1��&g�������U�2~$���-��' F׭�;��5t�-�\*_��aTU	C��i�U�Ջ��l��\imdr��ɤ�X:�յ��,�Ԅ��Ꮞ�А���TTPPP�:�`���"�%��(������ �K��RI�]���T�*K���HkpY�9]`���^<��e�a)H��ڵy[Wy�W�ਝ�2k�$�\}��,2�UN ���j6%��"��<^5��M�����_���^5�1�5=��֦���a�D��J�����!P�ݦ�t��JuF=`*ά?Ʋ�I�W^&�g�
nU�j��!z*7~����[o� �%.r�Og˰T������f�����aH� � o���XA�����EZB�R�+>6d��,H�C�H����WX�oU���B5�`��9l�D�)��ꈬ�c(��g�Uo)XU���%
�![c}��	����d8������ X_͆bY�5�/>`�a�A�v�u�bd�k�,b�����ǹp�~ǐ܏��+����� �mrf�����GM%�'����FNKML<_��pZ�,R(��_�L8u.*У���lu��[`�OQY���ob�	|�e.�C5B��j���3TB�'p�:���I����ޙ�ĠP�_3t���a.CU���䝘��y�;�{_$J�9B+ɉ�D�d�4)�r�#�����O2ɸ;R�ޣ�����HiTk__D�|`��q��؜:��gf�$�_��bcc���m<J�Ii� 6�'��GO�b��+w ��i�j�{8��� vH1}���,��l*υ_�*��H�C��6o�E�5{�«P�<ׇ��z��5��1��r��9�|��A�C��9x���`��qQy>����c�z� r2�]�>
?*���{������Wg�p�<� 8%��WW[�!�~��Ye�,���t���]�͐/+��~��ܤ�qJ7��:�����9km=,��q�H��&o(�&2�=�-
d�P��PEVM([���87�'m� �YQD�^���(�c�u@�o����j���NU�m��>o���V; �%Sa�Y���"�m�WDy�$��/E���q�d��C5��3t���lD=��F� ��\F<�	���c�V&)l�Q��t�f�..��cK�]�&e|*�Ź|(�l�K?!����p[Nf�/����I�K��G�҈��;tv����PU���=
��FP�#�B�XM �����R013S�a�r�y$m�XD���{A���{�n�Q>�.�E/����=�G��*և���cR2�����Xoa
���d�&���}nS1��_Sޓ��)���jqPog������Żj.827�̦����1V���_����,D���O�������h�<����A�
B��5�*�����R^���<���b�'����L��u~����S�V����{�4�ʳ�XO��($��G/�d��j�N=]]Z�׋�x����]1�	�;>�%��q��~��z�E�R�K%R���@��na0�>�ph�l��ECJ0�\k����YOw�Ƞ��(!����뀛�Ȕz����UU�7W"{B��3_?(��NS$x��Ȝ����n�9��s2�c0�^����G)1J��~�I�+��3��� 4��cA-�5��Ҫ[�����Ȉ�r&�ծ5\����>��nk�F��*]�=�8��m�-�z!��x3j��>�H��[<�oz�=ӹ%�4�	��YF��J��I0�J����4����Io�R�͹7�b����5���K�[\�&���l����&���3�a̘y�XϽ��?����m�����~a���e���(�S����Z���C^^B����X>�z6\��.2@�������ˡ5i0��UB���yZk{ii��޽Fc�����k�����=��`[)��_�Bu�3|����{��TF�8��"��G����IfY׽X0�^�Oz�"��A���R-����U� ���$K*�"`NceD�׬��'��A��,+�������o�f�)E���(��0���(�t8HM!�d5A`�?�TףΜq'�&�<�����x�/^̘R���,A�����/� �P2������:l�@Px��U�7��kD�� �9�"LFF!��
L���GY#s����Qx��؝����,k��C��������ԯ��EPƗ�a�ا�
�7'�!�o��:�@:�����ֱ���Q���"�k��]R} �?0�XʏY��M����]�(��4(?
W�)��8��s���l��>�6j��1�|��Q~N2�#���
��oYr����1�h�n��o�;P>�u�l(��K/���*�%˼����w}���3�����B��ƅ��ŠC~��ϙ�3�%ݳ��=,�e�y?��23����æ,����B��]�����q���-����<tX�ݟ�ܜ�5��X��ғ�n{&�9�J�kE��#��Gv��5�$���]�ڐx�Df��T��H��E�� G$�9#�ǟ�9B�4(�Mx ���=9 �el�A��3�,�5�[�ƋT9�8�ωb�A{ƣ�p���r	K�	���d� ����<�)S�A�=�(�����ww�\������M��Q@�������p
���z'�\L՛.��j�'�7c;�o����x.�W��M������Qh=����(�
E��=3;�@�@�҆S��tH�,��zt/���./BRW@���4�b�{�h�t�E�i��ں���!_G�۪���QdcA���.�����K橀�Kq,�z�D߅��p���R5�?���ѡS'%�mPEi	H��΄�X���UwE�h�����(;��1�k��W`�� ��6E�S �_�a�𶕕�/E�R��9j��F9��W�NF�Т��ĝ�SXPmuj�z�fu���|h�A�,�0 3O�Aˤg���E3j�RP��|?k��c�l��0��?B���*T>��Rl��O�
��0�B-�:��R`���`CH��/ 5��� �_�0�{܉��'i����*A����!*��׹%];[Y1��j֬�}�W_|���r����J�ߞ���U�0�.�~��i�'t��R�.�߇3���N��eF��~���ߕ��]\\��{`I���+S-��Ze��Q^��*Q�Д���������󣧑��'���[r�??�����܎#LG,�\4(�UPߗ��D�d�_�Zv�=����ߪ�&�E>�*|:�>�]##qԊ�����@o_���A��]�CU��;Q�{p��N���U�b��!�a�x�!'e!P����j�w gD�y{�K,J�c�>v���|Li��$@r�� 	��0������j��i<�~�/�H~z��cO{�e�SV��ڊţG��,��w>����)U�ub��.EX�*  ��r͐Jqq��qOڿ�ܟ	�`F�\�(1�z��Ш@���^�e�FfcԏRs��{k�4�tH���X Ex��s�<��g8���#�mٝ�5z�����κm�t��h#�{�G�\�YC؞'^>l�≮TO��GYHZ7DK8P�z-�X2�H�Y��Bsz��%�/KS�J� ��	��%���9�&��&*c|���d��I���	B����a�㏔gC�<��Ŝ'��#E�����ߖҚѡ׌C-���.�/,��]b��El�a���X-k��|��E��准��F}� �����|��)|�Q�9J�:�Z����	?7���_�<-ؼ<� �3
\�¤�(�R����z��)J66�*�$�B����:�+E(ND��~*w�p�hw	�s�YYY�c$�r��p n�Q9Qɪ13x>����/���M??=-vȮ���ҵ1|F%!Q1�~f��<�cs���{IU����������S�a*#�������ݖqP�+VV�~c5a����BHF��t���T�h�����M��!@`'���J�EZ��Զs���A�S(���\��@
�6���:e��{�\כ�����4{��(�W����z[0����O�f-���Ͻ��o�c]a�F����FiM�PC��\q;R0t�_fG|�G>X�g7�YڔL�Q�5����-�
⇨�d#�Q�^��4Uy�I�n��EH%�!G�������,�����A��X�SA%��7w��iԙ?�v5�4�9~5q�ᗒA�˷�.�R$E�'��/b]��%��P�lVY�� *�o���(Q,>A%FR��
�_T<�}�woqT�%�[�Ѣv7�GgҳU)����՚�2��<c�6Ӆ���\��So�jRW:��L���6�	�:�v#R�J������^k�F ���z����	>o5�2uhȾA�����rH���	V���\ɧ�X�c����30a;�4�3�
Q�����$;�O��e��y�F��I��W7)	E'l>�� �H��yR=psdH����:�(�G����X���K��Y�.CN}�O�t�������4���C�;sSYY�P<��Og���4�v�����i���tJvv6\&�Au�x` H'���Tg~}07����\�+SP���q�R]E� ���l�4��Vr�w�dU��
�j"E�Hs����|�:�\<KE&���uP�#O͓�_A�Q`w� 7"�����w�3�Pt��CQ�r��%0��p��ӣX�<u�ʲ�{ (�|~�(n���7�5�I�W�x�d����`'^���SL�; �8�����`�~ԍA��&�R�G�n�Q�`x=J���O�Q�o� ���ܜ�X�9��AP��'[�uETVV�6j�T)۬�XԮ}��7��q�;��k=FqI���9�k���s�HZ���tn���%mF\}�B�e�XO�d7M�vf�@1�s=`�{��0k����i�4��Z��/��m�ü(*����o�q�$O ŀ�uϷ����k1�s��۔��2�����5���>��3l%c�,��A�(��O&�� � V�.O5�@M�PH.�ȿ��KKς�ZP,G����gnc0�LoyP9�잫m�Oj�똩��dL�dk&*�]���.�î���*[I��"3��KU���2U����&W���?���³���@�sa�����/QV�:i�$&&F�LZɳ��-"J�"S0K�U� �l���ݪWt��*��ńب���ӌ�˷��\���^o�0,�R����,<;���ТH@�����)|���H~�YJP��(b��AZ�PF])�8���T���yP"% ��Z����<� ���O�����w�>�6{�Q��`ѝ�SBZ� ��ٽlØ�����` 3��HZ' |��?(��-�(�mCLHa��,Z�Pm�����~ %@GJd�96j�@{��OHJ���2�~�)�m�AJGD~T�����)s���3u��_+��h���j����g�OO_��ͯd�8�0�YD�Uf*^�;,,�cVo�r���k��p��xm8�9*�y���Ȧ*\�HA�O����"A�����7;Jt��x��f��kRaD�{�Oܸ_��)�E�<�e�U���]Ȉ��3t��N����Ap�)�z�yKlt���o��Lx�H']c� UK
�X1wMG�pBn�n;}�=Qh�6n4U���,�y�O6��	'P\�W��6���T���s]��!� {� ��G1W���?�T�з�$������g���R�h����v���M�2g��e�b`]uT�44�k��n����sU�z�O;�Q�j���If��7x�S Mڗj6]l7g:V:�W|q����9�Vk����u?�EZr$ګ\�2w/�lNF	��N{,����YՠYr6#��qMXB�Ѯ����1Z=m�b�#���5'�Q��"������\n������Q�,D�r���٪Kp�~�E*�^ۚ�L��6? ����ܘ�3�5���Li���5Ww6�����Œ���)�����\��ׄ���Z�  :3�}�97��ڒt>��ñp6��R1f�W=�_��?dq�Zq�;"��d,L���v�s$<g$����-����k[�cJu��Eox 0#�����R��l�;��AO���˼ �����j`%'/��'�j��zl����$�{}�G�m��z��J�?x,�q@�>�%i:6;O'&>[hƢ����4ҩ�2]����Q��@�M-�&��Ѹ!�@~�~���ux�����7<�ڼ/�M�^�d�pK#lx�h�WϞ%	G�|�b�X����|�摈���ę��L�/��}�z=(�V��״� ��+|\�]�J�
�?�K���O~�b�⢒��'���z	J��4ںW\�sd���6�W8% �҂U���O݅@�Dt5�2�R��Q�d_5Pg�O�4�a_]b�J�� ]�]��>���$����qi�=Ù3"�ԝ6�㍭Q��L���?�Cs�a�N�����v	E�@�^n�����1�m���W��o���w$S��]L����H&���^d-%'$	[�i�m��R�RQ&S�Sx��	�ⷓ�����%B�S��u�����hx�n����ka?F���UI?��R��\�Lk��7w����]_NAAݿ�c��e�H	��&G�O	(�_��Xٚ/Q*��+d�v{8�ͣi����[GG�U+W[I��fm"���ֶw�x��m^�0�A�hs���Ê0fgn��<X�J��В���Xyg;���f$�������Z��g��m����(�!l=��x~y�(@�ZIw�@��]�o��� X4�S�b�f{ܗ��=��[�ن)̶������w��Q�0�4�w�칞��G��� ����1[a���v	Lf^�p�)�y�MC��jU��Z�F+��=�'�=��!���{
�G�,~>��7�#���'��dt�7J\�*?n�R'x��kC��Au>����]��nD��you�4�������;S_~���^:������ޚ�㘫��p��H�[5�܄�G0aɱ8Al����y��}�[����7��y�
L�{x__	��SԶ��G�����C޴G���y��I��-r�'��CT�Lh	��d}镟���,khI�A�RZ�x5oɸ�F4@h� ������5k�@
�幱�pV�����+u$��s?��!6 ;�?�%6�S'
��9��%Gc��~�<����E*�~�:��Y��qw���[[9��x����d��Ȣ��� �U�L֍�&�A����W׿��7����QX!hW�9�4���]��L5Y�+��u�hј��9�j�����l��rL�K�pM@�Bu�K�����?ϻjc�����w2�� <���� Bpq��?�����=��
棟r��,��o�1�c�>�<~3С�GV�=F8��
.
���Sٛ+�[E�潗�\i�9"{�q�%f�I����Y�d�j��0^d���q�}(�cxu@�qJ@7d�r��I"�S�]+�y㻷��.+"u�ƞ�scgv�Urv�G��Go5L��F��L�Xb���Jh�)y�m��[p��������PՏ|h�Q�q�U��]��	��f�;M�d.5�uSY�N:$8� ��+�rQ�7�4_4ϲ ���
3ƞ޹1{`�N�Y��հ ��q3����۹�W�n?,O�
(�� ;Y�NX��J&]bu�~ U���Q#=Y�� ��O��~��#�M�!��H�E9˃D�"���$l�8�Q (�((��/���w�+����A�%"��_:����DlϬ��3�x�*+�������}�^x~$�m��S�Ԋ��aCI�?o�>��Ӳ�����g��yexl&��=�����!{@YQj�pn��*�s�2g���~����B���y��#E�ځ����g��Ybǽ{�V5ё�a���N|=;�.�0%n�V ��.5�ɸ<D�hP���,�$l'���rXF6n"�@R��#��ִ�E?�H�S1�kӍ�2�f\�rn�㡵��/�$����㿲6������hK&�o:����=o$���ad�2i���Ea���R��Ip���U)dk$ȗs���M�\ƣ�&}�p?���$��rE��UX]=i�0i�[�����	SR-��d��o�?�WLHN��'��e����R��<��Q�: �;���'���n�'�oO��_P�#���JG�S�8e¨�'l��D:���r�zޖ���t��K���;hH�J)�;�isl��/�h�4�*
��)q�$��{5���d��:�S�(�>6e���I9Q[�v$�4�-��~�
um�ܘ��fP��`����j^>j����$���Z9X1Ghgװ��ܝ�'ߓL���Ͽ�,&���H��@��fk�eO{l<�I���ܧZ��zntW��z$DL\�߽Y�&o�Xi�YQ(c���O)�ү�:�T�\4���u�dq����.�>R�P<��J��3daGn�A����U����,`:Tt�j9�dO����ډw��H�(s�ec, �A�9�H��$�!��c�ޚOE`��`��o�߹��i�ۂ'�REa�4P^���#l�<�`?i��~sE��0�bL�H���vGH�~̎m#�!���D�̱
h4�r{h��˳�5=\�s���q|F�J�M�Z�y��4���i(��V(�à���\��{-��rG`��d�Q�\4	�r��]��O��J5,R&�m"]4�����z�Ude��=��
�}�������%P�U��Z��c���܀�~  @x%gWI��!�6�KGW�n{a� G���~�+�+�#;�.����M��)?m�����.ƴ�)t�nZ
j�!l��OX���Y1�6r�P��-!l��ߓk3T
�dH ŭ?�M]�'��.��4(�S-{�燌
1,oM����ѓ���~N$����	}���Sq��!���-qĖL��L>�x�o�Vc�1o����Gc�i)���Eĵ�֔���?K��$
=�}Ѯ�d�fV�kS��ˬ5�l��h>�v�bx'�%��∠Դ��:叞 ��'jb��[8��&<��������$]���`��Im`S��RJ���&�����ޚ+��e�r���B��~���
C���w,N^�?�XB7��r|����[q��I֝�D��}f�um�d���8����)k��L��
��4���A�4���������&
�Vl���HS׽c��@r�]�8o+�S�m�]����5_?�ȼ�#��Th����,�P��M���������B�^Oa��E��Z�p����;��l)�K���$vj�'2R��B�ffkZ}�36���5x�7}�ng��o��uީ��qB�f�E��}��0�|�e�R��`k�~A�{�!\�es*.���K^�Ʃ���D;zQ�ՙW�R�X�`x _.S_��d�Sf;@n7`p����D�K�a���Z�i�нZy學'y{�,�!=��6���^�/�pT�ҙ��>qm/����^h��dU=�5Y?t��"iֽ��8�����;�-�u#[ǩU�7;��CRXם�N�.�C�t{5��T������m�wWL�RP�p9�l�Rj�6H.�nd�>�s�kRo��PRaf}��Py�Ɨ�^�
�bz�.����zK�	�����:�ͦ�2�0�0y?���r�y �(Z�hXes�or��V=�D�7�Q�Ƀ�m��ŵ��!
<�&}%Hv��'6`=�F�����؇�7�ou��s�9b+:S���k`����L%��`]�����g��[q�,F��iqGE���&��=���U�Zv[ge5ׄ��|>Y
����;f���:J�
#;�A���5� Ѯ�0����2v;�;�O1�j�kEw���X+kۦ �ݱ����]
�,o;F�ݵZD*_��Y�#=�nIs'�Ul������J\*�!j2�Hs�F�8L�5�8X}'�D)M�\�~�{��0)��j�)�?W�����ӣ��P����t/zw �\^�53��ibC*��L�4��YíRV����:����]{�(q��`�x+NV��(�ÛA�!�ɰԱ2�GU�ub|��<�>�P�W�VB1�DcL�uwԵZm7�?���57�.�ВYy-�1�j���.�,�q��H�b���$���*w��Cd?��{B���� {&��5����sV��y��3B�Wb�2/͋@� 7�	`�Zs��
�9$�rj��x�P�!�B��Cp��\���Þ,�Vy9f����p����LN@�Mxm��9��]��G#�L�b���
��Wqw��v	+��؝�O�=,H�.���3��������DN�?���͐�}gD���*�ĠS�=��\�i�\�ݜ��ql_��|�2I�[<�|4w[v��+��先�>k1ޛ��#c�b�x:�+++a��q�{J�P�k�{����Ѷ.\��v���=��u�.%�@�����/;���}d���!��E�Ё �qW-��&�´�3�n�k����˫jS����Gz���ǻ�Mx-�R��&�S�ʜQ�L]�)έc$y��9��%H���4#�[d"ѻ�����dmX����ՅY�����'^���T,����Ș�I0E*-�*���(��ɜ:�$��xc��t�%8��(��3g"��\��ze��`l���h	5�&�P(���I��^����3.����y�j:k�j� �� 0�C�?޽�P:�t���o��3�Vm۹��D���;����ց=�/$U>T�<�^���!��x��h���k�pX�Z[#�:l�$�a��~�ɽ!���x@��H/�05���\��K��O�AZk�@�K�1~������'��.��9�v��͍K�q<��VR�5f ��2�ϙ���/D��-Q'��j�s�w��N������Wk�J�ꗠ+�/X�l�]r��ǣ~�;� ʡY�^�*f3x�<B�� ��]��FKs���/�����	��buɚZ-��J�$�
j�݆�I�On+��Q:�:���H�k�3B3���x���$_����E��%�����w��ѓ�o�!��_�Y��N�+	���x����kR�	��p�X�_p�c�Q\��G�$ ����t��A��7q�r�������ϼ�r��.�PĨ�Ʀ���� �g���2S
�"zm���5؇� \���V����r)�y��l1�28��;(��oZw�]�=Sf�bWc����ч©h������T�,��������x�?���a7P] ���l榌��	ۡ�$!E4����m���7ي�v"Ċ�Е��p�3�8�.a����^t��û�H�	�!zqR�a$(�d4���t��{��=�� a��amjd<g:�<�!���	E�!�;���[� ������C�k%�-�N��0Q����b�[<	��\��9Y���z�b?�Ԛ��8C �yy&/��ݜ������wJ}"�T��RLk�?W��d+���_�ֵ)�@##��|
xk���$��Ճ�� �j;mcC� ��Ҥ���A̩S�����z�@��� �_�(�=�P�o�� ؝���7�pl�t��Lx��F��i���/��w-d���j�+㗬��y #��)���~�V���6��P��|bݩ}5��sL>��sB����ׯ��+��1[J��ό����b�F����p�r"��������0��I+?xRL��Ghh�Р� �����ZT�J9~d���Q̭ɜJ
�^�E�ze�H�52J�R��=-��N9)�pY�G�Ĺ���k�W�����~ǲ���
��i�y.#mw���&g+��yv�㇞��?��:kΉ�<=r(�@�7�.��~?�y��~��'����u�K���k��I��E����n��46n;�M�"�q�d����(�� ���!�,-��?�+���:Ny$H8L^��Z襱S}�}�!]L����?��IO͹x��_Ww������il�{�x��Ô�#��ލ?�'g��,�Mp'&��$���<�z�h�?iI��I��׾���1����ZR�<�������ٹ���I�Mh�F��b��?�S����.�k�ƌt$v�ի�������M������Λwn��V��쬽�J�)0�.t��G6��Fba����
�1�w�ڙ����7����˙FU��r�����ݝ�t������q����l�Z�����gP+�_��&T.�|{}�^zdf�{����������<���>��y�.u���b�e�C�GU�J��Ġ�5����ĭ��@�@�5�Y+��'�	iL:+.d���c"+�
�s��v�*}�ߌ�_�hc퐞e��\���N?��v�U2S&��zv�O��Z�wM�N����33a���b�#�����p��S�,�y:��w�6�pǡOnm�ɖ��m�$?9;��a���`��:�菊�M"@q$�	#���l����J�.����֚�ߺg��ϗ/
�����&}
d�2/;����.$Ȑf.�M��Ov�f����䵓����7�/1�G���}�{X��&�.�9q�!B���D�|���l7��mf���K*k=��]2��
;SĞ�/y?%�v[|w���e`]����ef����Δ����2]�v����D�/����G���
����G}x~/�Ʉ�-�e�܅{ZD��>K�99�s�"Wu������4��o+�Y9qsYF�r��	���߇����Գ��o|��&k�%.����L�GP��*5���&J�+�.g���'}<n� ��d�{�������>DM��������+j�R؊���Rxz�N����4E;y��]�h��4���Knp�ϫ|AaͲ���Buѧ ��W2��_��&�CC����x���X��� �o|X�����t���~�����:/���?���ǟ��rz��6�7ȡ�`vO�V�=<(�;����,BQ�I����c�ۄ2Q�-Ǥ�����A�]�~m5��->�]tQ�N<(�<iM �����>���Kn�&���7�k�p�YuIH��º�ѝ�;�D�-$W���a<\d���ӝ�F��bd+�5D���٪�? �=,C��V�뿴o�ş;[�f���~���0��׎[�詻o�ӻU�>nY�\����7��C�Ap*�Ҽ�z���qYR
����,������.jِ��>�bب����/�QGr��dTW�X�@*�s[���>~6�ꞗW�$�Ԫ�i��9���Z>�{sն�(O����Qk�'It�������(&��N���x/I2��+z��W�(�5������X|cW��d���E����{	��ӫ��j�K��Y����=>�#x��S����?��(Y��|Ztm��M�ZC�{�
����{m��%ټ��g���I�gp���G�Ô�k9��̢�/���m�o�.�ck�Q���S�9�E
/P�<@��Y�b����f%�)O0|,3Թ�幺�P�]�3zyͪg!Z�6N�~�9�|��r�\V`+���ƀ(���E�pْ̚M�����͝�y%�m�_^V���(/��^���������r{�@0���4\/ J�H�IJ(%1 ҍ4C����F��F�``�c��（��}��ﺼ'���g�s��ɷ��)�`m,�Z<SbH���NGAƄ^����(J(Vg
ƫ�-~~{}��f3��M6�V'VX��sI^�����]�� ����6�vc�e������B���U�V7
W�͹���n��j<bo���+�����]��s�LQj0g@��۶w���v�_AØJ5��P��E3TsKI��fbΖ݅���q�1jk���Q�w'ғF�O���F��]�bE��V�V�W���p�B�aە j�����3�3[�]�`��T_G�U>_r���Ch�2�
�r�� ka ��$W����n1�-�3ע��5��azO�!�Nl�(pD���ꊩ���(���V���乩��KN�iI�Qu.�m2�;�����U"8I��1.�
ef���
���|	���i��zg����c����g�����=�vvA�²˿�+�t߻�#P:J�f�����GV����i��$�qf��F+�1����M_�"�		�k�
	�e�*����}�x�3酘3(����u��1
���ٗ�'o#F�֜jA���,�ʷg�Җ9�X��~�y��^阘�2�s0���향�F�H������qڪ@��=M�A�.V�ƚ%�h�M���m(+$����ł-��a�+�~���I�/�X {�`y݈���e��n�5)�+��!66(*�Չ����5C�z6�W&��������ǝ1�����Z���;ga�d!b��-|_Zw)<�/�0}8o����O���g��B �AӪ��e��c=��5*v�w���=�,`���dw�D���&��w���IB,f��+�F����=��-�gM꼤�-�']��2����t=w�=֚�~|�^ �h[�O�x��)-�L�2�Y�I��7�¶�=�r�%�A�1M���}<��s���o��y�T4��LG�l,r���=��[�ݤ6�vvU�zs)��q���a��n�q*��!��@!J�y��Q˺�빏���'�K�iy��k��h�Q����H5F�m�$W�2��/�&'78q��@� ��欐��;������i �3u���R^�ln�DCk�߁�8#3�Ҳ �r�.��ӿ��&�M�Ò
v�A {`���1�=��n�k������"ٸĜ�[ �94af999Oј�.ѕ�T���#�k�X7��-^^��T�@�mM�!_|C.�ӛbL>	���b�k���e�$+����,� �L�ƶ�����-.Y�Ǔl�t���F�&i����$�D��o�ae(����}�k�Հ�����G���;��HF�#Q�	��D� ,K]�^�	*����3�Qc�׮�o-B&!�M�TIg����홷�Sq��	�"e٪Y^+����ߜH�z�Ե�c�/Q��d1�1��%���9n7��׍7Ϻ��	5�,OڒQW��T���@�P���+�h�I��F�GC>^N�'D(r> ��~���W���J�e�'B-`�7^؞�;�y��z���1���≬�{�4h�>&:K6��-����BII9�GKw�,�(�W�j0���C똨%rU��:�N0���ʹЍ9q"Ef0i���f �2,O�L
@v���o�*��)��������@�5�ݳN��
;DvQ�n艗
c١�*/���ؠs4�<ԈH.A$Aڗu���İ�+V#E�m�������D�1�A ,VD�϶�5BH��/�����!ێ��t�o,��ebio��og�Xi�(�*ǲ�ݩ:0�1�&Q���K���RW�ٷe�0O�7��,oGoF���[^ECiP�6�n�(��@��l_6��vֻ�x���?�T���`��ll��mj��FK�R.r�(ë�v�>�P$&&-�����S$��!L"�uk���֩Bx�+T�Mk��P5z0x��li7�o����_������V)�72��g�F�_P(t�$�q��ׄ��(���U������2n�z7Mr�j�-=q����&���G����ې[�|?dt��E
ԫ��7�B�`�i�2^���쁉�O�B�I��Nzj�8��/
qP�7� �>ו0Xd��M=����ݻ%NX�\�R���\E�`ࣕ��붤Ӭ��q�\�hd�|u�G��ʷ�r��*������?Q.��^a��gI,�o�9�"��*H<ƙM�罶���cPt	��<}n�X��!~m�������q�
�b�IJ��[<�|�Vm�>�b�
�����R�A�4�������]M��{gp��X�Bl�J��Y?�a���k2�D7�+����A��&�G��YcQ�x��o%�(Np��5k�q�ٵn;�]��Y깱Ч*+&�dzl����=�@M��Un� �\���mik4�f�~B�e��.��\�c'��&1������l$�N)g�
u@�&��+�-��#��Ltk����U0uJd��{J�;9X1�����ɳ>�� ?�R�.�ȗHZ�e�N"�Tbh��ea/�=�~ƈ�oj���z=��Z�&٤)q�;s��1�l�8!���Q�e� ď���O6�ժ�����k�����OD����W��-��9��@T	X����	�f��)̤*���������`���*a��h�����prGW�s3��;8�!}���HEdD����`g���	Ҧ?�߻�O�,�����޴����3�� /�$�J�e�r�_Fw�]mP���Sx- `���Y��Fy'r)[Yd�0ի<{��A�ɴ5�!��$����`��[�F;Z�R�ز��7�{W�P�$���ѝ(�Gְ� �����N/�}F�ݍ+���uY	����r�y�W_8TU��;^��v�!$��Do�)2����'��^���&�lW������3�����ޖ1,�~D���s�A�c���%�݃�b����LW�s��m�~��s3�f7�B��5��Ϟ=c��*57G�厖Z�;aGo����=�x��T�^�Y����� d�dϳ�������'���^��ʪ��8���B�Rwm��Z�h�[ւ��^)���#�#5?��Qْn�ޛyI�w��D���e5�E,�Ёa��ɖł�C�u�ˤh�R��~��9��Ui��C-��������(Qzל�a�t��Qifm�Z/�P�����e)�G�S�p6��р���mq�TTJ�q��Tî��d�v�e;.�fE�<�-�c��i=0�
�٢=�KNQq�+AT�ý�s�g��I(�THO���o�q}�-��t������h4�PR�0{rq���\j�/J��s��3c�\x�`�����5�h�=�QNݞI���L�ѸTy:=s�|8fa�z���Ҿ�I�a�ϰ�����@6��,*�NΞ`Q��)[KH ��R?|���jT�3N	�S�F��*��Z�mn:`���m��XT��zZz:
ʐ��Z?t��5�/\�}.1f��f��2���̑B��QV�t��gO��#oG��	�@it* ���*�S1�ތ|�Ci�E��:�\i�]a�j���g_�L�Aߖ��i���r-�ҵ�#�[��}C��`jC�cM��X�,h
qj)RA���o�]Ų	�8-�^I��ܛ)�&'�ՂM�"����i��G�����9�p�M��4��Z�CP 8;�U�[s8/�}��P��br����-w	4^���N� (Tl�"��E2�E�~)�i��T�T�
h�K��VBz�m��1��),�DYn>ⵉ�T��U~iz��� 9=3c�1�9Z�7�1������3|I�^M��|ZD�����W1� +"iu���L>d�]�����;��ls}���g�x)�_�\�7#]4��?��pn� Q�a�5�}՞��8�����fS����z���F��Jo5 �D��>s�Y�p�F��}��\���kD��,X�>�v�>�*|��S6m�f���tchK�	�g�㶽ܛ(�V�Ї9v55͸BA���+>���0�����+W�\���(,�a���M�v\������%���!:[b��8��Y���$�/2�us��W`�|['�v��D��ɳs�*�{�:Km�C8xn�>7N�ׁ�s]���� b͌d3����aH����������H�J;;�G5>R�^Ж�#������݌���B
�X�u��;>��� ��ծv^9�x�N����`E��NV�,,�C�:K#?oww�[�H\PPԀ���V���W�ϥ�������Y5�u>D�O*��E���#f.���j]���bpe�\Mϣf� �614���"*�=�b���qi��X��-�c`J�܄"(����d�o-d��A=��6)26.+6��[8[Ζ���u�8����t�ri��._�,U,��^܈�G'R���}X���N.��۲ׯ_�P��db���uiniaPW�VW����b��L+((�qD~�l>2{y�����p�Y\���	�

��җ�yff��z��*5$����=�%�'S�0Ηƞ��������2��)ZU��k��Bd>i�:�<���ǲ+��÷	�~�(���\� ����q�i��%�Ţ�3O�C3�Ԉ���b��MP�A&'V����Ǐ!j�?/��ʕ�7KI�������e�������ϊ{������w������>x-E&%�~MHy��Mnn%���j@��u���f��}ˏ5��+z���z񹄻t�$\X�����n�&�c��Z6����N�p�,a$p�d`�d�*��\�)l�Rq�Le_{�)�(��J���ښu#��O#�9rm�N�A�=k:Ԣy��w@6Η���n*��ώ(�~
�N�I��Jޔ��;�!��Д%��ţsi_~�>C]�� f�`i	�$�Q�9	�3B����.�K��*��
4�0y�ʫ��,����;�w�0�3w�k�V6"b�e��5� =���8���9�XG��T�H��±�d�t�}B�tS����`@�I5	�= �u�����x�� a����W�G4���G�G�9��fTI+h\�%w����i��%������ʩu.��M|!�N�k�3�۴)`��K��,��^�t»�����~唘{�_�b�RF���2F���S���EL�Å�%p����۰�<�n�1{�d�ڴ�A'͡ˌ���P��?�V�J�e�G�z�sz��X�m*�3)�e[�3�fh;��[?] ?/{>�F��pE�D���<�_�I�x���Γ \T���R��O��[ �a�i�<jm�	K��#E&:�H�.�ug� ]�{��?/�yb�L�WD���d�^r�
K��#Xg�Wll�0޻Mv��pG�_M�qZw��{���E�`��C��;yf�A�9�����Bm��X�[��s�H0���de�F�\��R_��\�i�Mf����䤠+����4�eg�fs0bm�GH>u7�"ހ����	�*�m[!"`5ʽ`ci2WV��A��x0��egP�	��t�{�"a�U�������~�2�[������|~��'��Z+<Ӕ�y+n�gd\�;�^K�u�a&�I��}�o���mԘ9�-��P�K�N�Ԅm�nL8�>��m�O�u��[���"]��-��*�iU�Z��?_^Z� d�-'~����G�-08Í�xK1{���^�>�i���Hn:���o	�~�XĿ{�=���#Y�W��Z>Ya��	o��b{K��\&�z�����f�{���[�BzG��*�O�֖�KE׮��2���Na٥���wT� K�N��l܁��1����-+Rc鏙��ۼ䣸���hc�b� �ETV~� ��@�1�}Y�~�P
�	e�d�eQ�[����U�5��jۭ6�j���<�c�(�)NAa=_`�Ym��2��HX�ڇ�:�5�r�{�T�5��)#;�o���:}��o������J��n���&8.2r�{�2��V�Y͖�v0E���g	vk���Ll��,t:��
|	�A����Fy������Wtw��:��T�v�������[ �آ��F�8h�d� @��B��]�K���[�
��6�������a�1��D�n������[������<W�,[��1`�	�����4�a�D���������ގ���M���(`�k����*���]����٩��G�3D)� ׼u��ھ�:��Y ��x	"p�f	���ES�S|S�4c�WN1�_r�];��X���^��q]�V��A�3����i1/?߽x7����6��cqv�1aKa9�X����a|�L�����RDct��L�oc#7);��R�H#t�+«� �������G�Fr:	�L��,��"�b�0/���i�)"��`���|l��� ��֞�&t���
�t�s�@�@�^�4�*�b��6���B�Bw*Ф�z>S��n*�y�[g��([��(ΕZ�LU�R��@���M�
�
$��D�%�) >]��π�����ek�b�SC�$�m{�H0�N'Xz3����9^���F|������3��{�B6����-��g4z�
z$�~��9��r���'v_8JҸ��c�]��9G�D�}�K0��5�}0O]J��9F$��N��@�M���Dtț?���������c���x�o�z��S���e�ZI�>�`���)%���ߣ�z5��l��U��%�i��: uf������ϑ�X��3�0�k�ZC���<<
õ���/�ϊ
f��Ǔ'�9�.�<���٣AX�k��S��" �Ǘ����x��Ps�m�?A8FGKd��H��9���J$\p6�c�Q�S�n�pF��j!��.3ǖ9Ů��ok�� حw`LIZo��6�]fU"��X�������m70�tw����\��uKL���%hD�kKVF��L8�p!��,�x��÷{�U�קo�ȋ����t���\�%�h�$8!J@E�>�9�?����������	��[�UӀ*ȑ�Z�R\�������@�0�yN����L�o�]��s����h<���݀wZ*��aMG��RA1�X���4@�*F#�a�EVT��]����.bR�z ���=4&r�b���"C[]qSBUig��t�2׼�Y��}["��fY%�����2>�(�ӰP�����]�I�S��1 �{����_J'=�Q�E��W�`l�c.t�R��f�|u�M�8�C�}�/�b��UH91d�P*X��CZ4>m������1��MaoG(\
�������]3�iȓx>��I�d����?M}�b�Ň��+�o�QN��4��8R�}���j�	]�]u��8B�_��4g� �B"h��m]:�J2��/ᰊ��N������><�W¬��ƺ�h�C	_��܉�)�D�$�&p'B����w:�/�S/�Qr�t�y�5�e���9}[]M����?YH��MtU�u���}�#�e'�.e?����]*�h�}8��h�{������ma��xr_��XvI��T�^ն����-e��m:5�0����b�d���3�JG������NS1x�m%����ۇ��q���UDJLyi�(��]%\)�RQw.���&�{^����A�6�d�����N�}?|�F��Rȣ_����"�� �\[��Y����uS��o��3[d���I�z��'꬧�>9��>b�k���{�
�o�a���`5�?�f�|��{(����0LC�?�@ٷ@ݤ�y�w���� 6)1���&4�Y3�tQw�}]�r���ӝ��]��1ټ]����TO��x��_���r(����7>l�B�1�7��S���� P�T�qc�m&��b�e�ρЖ�N�.YVGR�d�ޏ"�l|��V2��D�?:��8X�'�I;TsG&�Q+ڀ�|X�p��qm25��[U��B�?^'�b���KGR��"�/�������?�e��S��tv�B����^!��Z0t�͇���f>�q@���s��D��f�â^�3'gC5��RbB��-{'�K�lhoG�ڈ�����vwX�-�����i�ŽE�!@��,կt�����r�"E=7����,Ҵ�+��_��6A~�e*��m�Ş����K��B����]P{�A��vQd��B}2�W\���F�YP' �� k����r��ˎ��,���(��w�U,I,}U�����:�V�Wډ���\(��p�<�E>p�U��Hk�z�m���iB,����$x%�>Q�9�2��C������^���`p����ԽסּN���}�s)�k��~-�f���+ne����2/#�b� 	�o;"h���>��ww�;�j�}�X����pb<`l2C�;��ׁnI���'g.�EWN2����&�2Y�OZ�v��LTi�/�L=�f0�/�N���_�yT�$��<�T��/^Y%��>�ޫ�@Q�Mj�%ʒVE�H�������{�>H���1~W��r�!t�#V����x���QW�����nײ�*䜨�X��~YR��l��s����Q�J�v�������E���B���aX��%T��]�`��a	W�!0���H�
�2�J�{�%o���bq�II1�q���%wN+j~~mUO�uk1K#ȸE��`�6�d��4�(3����&��6/~0ٚd"h\_��gj享�'!=T�/{}B����Sm�z�V��]$ʾ�X\z�'��6f:�=��rZ�͏��n�̌���u�F/���fM�����H]�t���8h\W���v��Qx��	]Vt1��.�S�W�?}�%k��T��">̏o����Y��tf��G���@mNH�.uA�4pe�p�"����ؚ{��MN�&Qr�XMe�d��ZS0nu �O�7>.j�g�O(�SW4�����8���}���7���?����ZM��>gT�T����$�Y÷a�:�VTޒ4����?�h���� ?�0��c�����.N�����7��d���$����FYo�H��Mi�`��$��(��/	2���	��	v��6��CF�͠E�������+�� )V��Ft"^�Q
�dQ�ٳ�;��}-j8&)��wf*�ړd�%�|`�
k~��W�����B]���W�^�gs�Nw�qT<���Y6����`Cr,�*R�~���7ž�(��˥ļ��l��"����QW�QkV-��)}���eևoL�~��t��<�y��'V������`2&�Y�WH�><�WahKzut�������}��+�w;���
����7�d��l���ͬ�_�*�� 6�G3�E_��;�� nJ=�{;���R{�O�Ԟ��e��� xhuA�_r�=�&lg��BH���l�2��~%����U��:G�j]�V�y�#��pPx��:��L��0�k��Y�����"o�4T0�B��p�O�f�9��A_)^P�'��|C��j3Q�R�^~t>B��KKW��kk��7����t��
�H'<u�O葽8?�o����^�%�����������+����Tr�$2PҦ9[�HM|��0!..n^��ؑZOg��!t��X�:�,x�����.4�����F4J�L��I^R��"+�|t�|P����;�?������+Z{�Rʁ��z��� ��u�]̴����S94��d}��G�|^@��Z�,��D*O@�iS(i����Z�b����b_"�X]7z������ ǀ7�� ���!��a����n���6��)�fa��P� �F-��0�� �(ȵyY{�P��t�����Ag�~����w9�)�zP ��.�}3��Z_���U
;��~�9F[�DN4�f�VZVb��pJ@�~+9T�IKő�k�����nk͔�=]�k�����1���ڷ��=e�l�pVf�2��վ��%��#�d��$l�AM�d�y�
s�ni�}�l"��{�!�#�?����T�ǌ���[6��O�)����x�	W����;�҂��ŗ_�k��i���;(�.�9r�$]���Tv1�o+�4�����	͛���[����2pJ{q��|)ak���L���_�3����Q������Fba�#�	����@��q�4鋺 M'��>��n5`��oڟ�'�=3��Z�iM)߯I[�<�[��3zw�}�Jmb_�$S���G��(�� ?��n���٭#3a�.j�Iq�f�����Z��Qv�c�����571}�y���+�G�}������G�_vJ���t`�3��=���,�븩�T��	�6���������j��0�kރNz;�KE�L�+��v�1EG]i���tBW'	ʋCF%joѷ���pBk*&�|�8��kw%<�1�o��T��e�!L�B�{}�E��S��4CJ����N���t�f0�e/�/̿j���Tu~�� �!'w�iPq�ΪR�>l|`I�}q�5Y��k�Z�+9r���;$�б6�� s;���W���C�H�xX�i�z�?�ß<|��-���� D#�\�#��b�׻Fq-E7���) �4]�Lq��6�V�j�2�苎�c�=���ajҀ�`�˘�0�+z*�X_x�r���8i���D��L�:a���K�H�_v���0�&���Pe::�-�Dv,i���XS89�6���(�@oz�#�MNT��� :�p�'A��B�"���rϯ����>��3{��s���z���x��޾�T�֭��0_rF�PIdqtW?�|�r�R|��`���r��%�		�<�eCDƩ3i�nܐ Q=�1=-õ��\yc��Wl���&�;� E��ܬ���5%?Y�G&�-�X3q_|{�5p��-���1�����xN�?��Mx�8ƥ�L�
;TG��w�ح�պMU/�&�����v�Xxh%Z��D�|�;��x�i\r�%Jp��b�l������{S���1����K�V�r�8�D�Ƌ��������4�&�7�77z���W��`	��@I���.��n�ΚhK���q��r�P��5F�̳Ӝ����͔�/nv�t�M� 1��Ր��S�Д���������-��3tŦ��#�2ےǛ���m~��D{���li��6}{�j��w_������!$�a�nl��w)��oD�	�����!��m���7�b�?��yk��ф�o�(�.3�P%�����-�փo=�m����2�	��9��t�H�x1Q��`ŨNg�Dj�'����n%^7h:���R��ի�?��K>�M�@��o�黼�M��@ul��<�zu����Oo���2������YRP�r
�^3�gS;yiIH�.�r��3�YTϏ�C�y�?���238���^������ÄyZ��)1PO�O�3Q9����g�EDZu-[�Q�c�� 21ɺ�wiltV]�!���OO���J�,��,s���~|�qü����O�֗�J��8W�&��<�5A���V$�JvS����������k?Z(�M0�D���)N�Y o⿶�<�F�|y��={�`��F�H���Q�-.�|���[0ўG��$��~���nӣ���m��� /�<�p��ZJd��r�P~��D��MDml��00���z��7K�M�,̫a0�g��e�g���8C���
i��v��v"���;����;_�\⏚Q"r�M*�#�r��b��M�Ck�'���t�̿��A�%�r�'�A�w�3bR��>���֏�U��1�
(l;`�����0o�1YF+���K<�B�`��1߰w��%�A;�����w+����F�\[�A�A��6ůE{�7����q+%�oT@qt��9i����"s�B<rL�YU�'����~�}|?gښ�\�_�ȌPqH���qqw:/_�o���+\��D�!��x:������髳�J��̚���6��)1��^WNk��$m�m��6j���4 �U�jz���U�k|�X=�A����&p�3��E+�����(��(<�հt�kD��I��&�x���_bh�xY��A8�q��텑�2����\F�jDK����cʹ(>��M���ny*��
T�JO�Քގ�?��@3�[F>']s��b$�(������W���l}N���kFl�r��H�i���Rsoܩ�/�_�p/?EQ�h���u7lJ�՗8�U�Nx�ME!��ξ�@�9��vZ(��@/�,GC�iw�%%��ĦS`��@�����j}������˃��˲��p��z-X=�ҫ+�7���')Yi�������KU����<�j@��sh1�=:烥r/�u�$2|*��{{�U�W�ܕ:���I�{�C�:�d:?ç�J����r�N4�3��ɑ;�~w�a���]n���{�����_�W�i�/LTu��
]��*)�O$jt �*^�~9z���� z�pi7:�S\��7F�6�s�}�yf�NCzG�v� ��Kf4.��o��rF��j+\���{l�'nQ�p�l���s-,u���o�9�������\�>H�,��2s�� oTK�Ԛ�߫�*�j�!rӭ��h,/�SF^] ZlaOR܆�X�cU2��@,|�맟��il� ���9P��݀�-��r"�ׂT �E�,��G?nw�'����r���z��C��>�h�p�nR�1%4E����b�ʮ�����~�Y�{&6�fkFy\
̼���ĥ21���߽ *v���M{��>v���a6j�:��e�P'��6b���}H�A��v@���wlw�����S�')�[��R�9�Pl�n��-t>b�P�{n�z)C� 2g�Bq�
��AX�����L�0t�[W�?��s�kYU�FWUثa���ʵǃ򠶕��m<@Z��qF���gr��ط��9X���w-m-�p3����?v�e��w�R�/�l��ӛ���ތP��k��,��F;?*�;��᧎�^�Y�h�z�%%�����HT,C�&���3<`�]�^A��qqP��9�9=���wbӵ������qX!���ng�o*B4�m�\o���S �%�I��>y�Id�p*4hq�8������t��zܖ�z]�+ɩ��&ѣ%ɍ�����rS=���������DA�G�����*|�]���+:��~����(	1
�K �ȶm3��BO0��iY@�鋲@��?�kb����!���j�ԵK�z�^M�:y�iX��L u�fM�YC�]��h��	D��c��s�?��S�E��Uȕ��Xx�S�h&Ȗ�˚{�{�8���<}��z�0Ǖ,�߀Ts}uuC^	|�'�ﶅ]���G�mk�BZU��w���K �7M��N���ӧ�v�e��i��ǒ���8�<D������e�6	�@(;�͔�ޥ��@�A�����>��Ta�ʺOAR~q��8��ߛ�S��[�'?�
�(�o��$��,Y��1�sW�P������@�J��F�[x1���Qr����#��쐐pPl�znΌ��p�ۡc��9����A�oh�<8�_t�Ǘ�٢w.[��W��O
��4�,��jT����ʌ��W�KS�4�����UB��}X����j^�c0{��.�'=t;�ݸ���Uy�Wm��ጏ�[�q9�,Ȱ��0\�MK3���Y�n����_	�&��Aסs�pm[�Z�>f^���T�y�q��q�ߺ/��^�#sE���l����F�Wq�{����qz�=d��(/B��	BH �!!�?r�K�����BQŞMa��|
tW�V���)���hP~�ZF��޵�{4.��s�p�:.�a׏D���|'�r��>�/���y��$tm�����lx�M�Se�v;�Y���L}mko:�c�akz���d�3�q�Kd��q_CL�,L��}aL��O�3?����"؝�┲cʤG���}B��W��I;�~�|��%���ܟ�����D�"��@.�c�%���o�<{�;�Ʌ�ݬ�5R3��4��6���A����
�!S.�Y��67�o2����X5_��t.ne�U#��%��h��݄<�F�Z��j]���*��=M�-&��:(h6�����}M�>}�r 1ǵ�$?b�}�>��v X�֢��|"�s��J���K��0�8\�v$#��N�%�?�{xT녙�Ŗ�I����,E)�}�צBo4�'�Mz�DN�b����W�m�S�k�C�<9�|�'�mizs�=�8�'��kq��d��~އ����,'�����z:�r~��i�l����$
�ZY�RL�]���A蚹�nv`WY�~o�&��1Q���!ç��1��#c�Ti��	�$j��X��:C�l�$�J���g�'M�:���KJR|���8�ɰ�ў���c^�)�J�s���4��
��~J�;ہ�㠱6F�D+E�;�/c0ɹ�w�p��9S{q�`�?�:z��d4h|iq�|����=&�z�+㯞N�<�ZH���r������V���[��M�h��V��f�ˮ�)Q+��2=5/e����#�f�"C}�KXNI��^����RV<Y��F�X�)%߮ć�`
�6/�;��6=�}\�}�/#�@X��1���0KM�O�"��˿�#��p�8�*�YV*C�U�Q��T���PQ��N~I����ug�%E0�^H���.�7N�_�ޒL�J��6۞����C��C�8˙�Ƞ�Q��q�j��4vt8�ԃ����A!Q�r��S/O���ђ�{-@?��R?�s�G�s�6�A>�[`}�%����,?� �yopC�)[�o��Š<*>4�E�����\�ABI[��_�-��?��9�������C!�/E��9�7|�[s��r�t�ol%Ք-��X3��>]�-vX�|����lI?h\���ՠܴ�uG����j�c@����|g�JME�[���m�ڦm�=��8Z��$Cx8i<���/����C�nz�v�M�{�j�����D(����zf��:+�g]׶�仓���9}��!E�)vG�ڵ�E�y��{Ʒ�z�b�w�пs��[lqEe��l��zM������s��5�	[�9R+<�K9�3人�Hj��X��z_K�I�|���v(��F�\:�a�>�)z�E�I$m�4ş1b+m���c�B\0���)s�N�$s��d��������1���c�m(�(�c
�8@�gu=������Z��HX�4��,*Ҧ�&}ﭢ\�X:�Wz5|(6��,v4��a��E:����L<�st�j��_����"���joi�.����̨�ň�q��8�1ts��}�{S�����/��-uw�ئ�$�,�׊�+h*�զ.D�}����|�!V��/F�*�owG���L�7�Պ[u�H���xU�0}�y�@s�����b6Wx��m��D;9!Z�Hv�-����xϏ6��AM��=b�t�`%<���vV�
��y]���y61V�L�Ue�Ig�p�����R���UT����JG{�2�A��W;�k��!1�U��Ȥ�4���t�հ:���h����t�m=Z�U��PFW���2l�@Qx""�����\�
�j�u���%��z!�H|��%ږY�hT�YO��"�c�����K#N�ʂ0����ݒ>PlK|ZCa�ӌ�g��p7��8����=��z|Ɋ��K����7wK�#��#��Zǵ��+>��ǫ5~��9qr��"�ɀ���m��X&cg��yM��7��g"�9��"*��a��	����u�/���I�j��Z֐N/�)'F�����bS>�}�]�1fgY���
�Z�^�$��������FMY�!7<������I�j1rzI��H �P�����K}F�:�ڴ�؏�S4{��u��J��9B�[ҭ9ŉ����o�ywW����'��1�P�Ӻ2&�Mqݤh��gowRn�w�`���f���+��2��h\�.�5:�YP�Q+R��A �Or�_��G���]�����!����9�:�L�(�����z��g1��W��֏���Rڕ�;��@�i"���cU<�:���o'�i�5�|?�����¤��-,��J��r���H��36�7��]u�[�4��W�Wk!U
��Q����d�f�9�/q���雗L�B�W��ύш�����ڬ��m}O网�����|#PrֻC��4qVG�[jh�K��n��Κ���2�Q���D�Hy��t]�,0�$�P��-@����=0�?pYEy�(߯d���+w���ф>�T<�◽��u�-ޜz�5?��̠��� �Bv!��J-��ba�	z��|����7e&�&� 2@�\��&�z�6���h�#{�A�ƪ��˫s�7��ժܯ�ځ؏N|Z��>C<������ى��ڼj���a~Q*+�d���0�>ӓ���SA�Mol�j�s��b1���9%���+EZ��ᓒ2t8�AW���R���Vc����f��3����]�j0Hx�P���3��6YXI�d[ۂ����B`��{2)�M�"}3��q��5�������^��]]��Ơ���L��`K�i�J|Z���
�IUOO�x��+��d�9�P�	�ȥ����a�@ϓ̋�J�>_�~:hI�N�]6]���Ǜ��Jft�]���/�Y��*��gPs���q$C��)rwnq���mo׽-�����\�R�������l=MO�����&{XEN_�u���5��>)�3z�m�!:Or[�܉	)��^����������I ٍGF�HsnM�����c�v��.g��0�Z9�_c�L$L�'��ozz�Gt�!iz����U�����u�v��it69Z΁з�~�ܖd�H~�p�1&-��#o�������pV�VK����}�I��9B��s?.�$�5�~|Ë� %]=n����,Ny�BEW#L%,�K���3�}I_�'�7�A�r�7�n/",�ڋ�;����J�q������Pl8�S��ti��/̦�Qmq�������b��@��Wk=j��<0?>a$� ��l�SӂIЉ�S^�P�ñ�C	y}�6ڝS��ׯ9L��Uη�;������'�}��je�����^�F�o~���Ɨ��k2���㓴�u�]}�x���\�C�U�u�B����ޢqޫ��_֬�6Z��SB���6���8��L��*,>�)�x+��X*¤����+�v�ߤ�]�5�����b;�)R:ޜ�����7��Ж�n�st9[$�5��o�X��q6	�n�C���mLw%=��1�����k;ﶛ��bi�,�q�!d��K�b�9��c�EX�sĹ��a��d\��B�A�v�'��ۨ�8�����3y��]��%���<~�>q5����|�~
��z/���a���N坹1�bb3�+��;��$r�ü)�}�k�:�^�Ui���`W<��JƆ�!���eg��^`$���nJEpv�-�{�~E�F�fA�A{a2PƏ�c���,�0�y�������뿕L����!�	�]h���2GJ9cBh��q��vT�N��f^�G^����Q^���tީ4WC4��!L_d���S[��Q�5E�Ɛ�	�A��Į��fC
�@>Ar$-����k�Z�����������%�l1��1b:,�`G�DPB	M��G�g�h��"�hE�QD2B�-J���PS �H��@7�ؿ�~`g�Ý���=�=g���ǿ�r��f$�R�)�@�v�ޚ!U���i~�e��Xà���s�Bn-��[!Hm75�.%Δ�O����&.�g}�Ao�����c�h�B���8c$,O�	>��r��4 <� �G�Y,)J�#��bx����&�(�����]D�����ew͹@�7��%�cg@��H^")m�veݻ�a�l0G#��e�䧟 Kf�Wg���rI�bKu!�U�Î2�m���4:+=��cOB�)�����?����h�[bQ��"��93�ui�S�
�:;C��UȨ��JZ�<%MAs��l/3�=U�	��ޞ{��aድ8ҿ}��H�T-��%�3���)��~��q�th�pC�4��/R�{~y�$z�A����א�X6S�1	JH�mb��v4S�tn�x>cZ��(U��4>�����n��}�DQ���D��L���=�Xm�^G��=b��7$N;����,���G�ҫP��J�`'/�����I��N�/|��]]o�(DE�h��*��P�А���B��/�~��Le��YD�Jv�?<Gs�)�M�o ��`Ks��x ��7��:���;��˚QP`%�22���������|�r���S��4*T�Y����ktP��Y�j��X�=�"���A���CJ���:��H�!�Sn?*��?�`�F�|�tr����c*w0�*_B��A��ۃ����/����ö��nHP�:�J@n����v�y�b4]�w�٦pql*8
����U9��9��s�R�[{���;����a'���@�c��A�Q�AE~�?@++�õ�)G����f��2�k0�ԃ_NCvA��c����<�-K�D�N�bl1�=O��������MI�6q[чvU ��Q2<�!�r� �������(�&�����G���=�"�V��AԪR�H��w�ʦ(H)TD�/����̀8r�f(��'��P�e�ygl������xqLH�u��σ�lչ`{;70�h��
�T_��M���o���<n���JW�����1����S�5�R<�}�%�[�C}�c��]z؆��ٖ���nmF޲Yodp�^lX�ϕOۍ����^�L�d�[oi3,^1���˾N\�M �f~�����WLۍM@��Ts{�ϥ:Y���dP:�����\�Rl�ѧJ��+D���5F�` \_���+�F@��y��c�TWw���'�������W2��ywA�����mof���@�\�kAm������� �l"^l����=t�5k���JV�^4�,�!s�9�q���%��� ���Y�Onq�6�9�d��"��'+YC5����[�u�_PK   �yDY�TV�w'  r'  /   images/3b67e01d-51b5-44ff-99f9-fc90dd618da0.pngr'�؉PNG

   IHDR   d   �   ��]s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  &�IDATx��}|�U��3�$!!��BhBD���4Eѵ��kw���ؾ]����~WV�?`G@���� �#�$�@B
��>����M�'�@F7���of�y��}����s�/�
�7dE�50���3C,*����*�@gC��iK����3�?.S9]�b���� ���-���-�|��Qew-м����`AUU�cGuך�cg�|J��*�Q9n;�k���*/T9����T������ł����V�ܒ\Y�Pn+��X`����)���&1H�NA���]��6�m����y���뎬�{Gv�=�{p"���D��W�3�">%�Uv�Lf�c/Q95���Un�82���Sy�ʧ��G���Ǚ�U;wi�ӯ��C��t�i���E<=�ibƦ����0}�t��ԫ���o#-7�(�|R���T�j�4|O-��?\�G,:�C�^��'"��~������Š����C���'��EO�mӶ�y$�G�GRVVZ�������Iflw��Tm<A�P8�2�a��#3�Q��)�ҷ���/%U@z��]�Ƣ}��6��0�u���Å��#k�0g�9gH�J�TRC!�6t8����v*��ƈ�Fl�\�fE�ʶHޒ����p�4��s�Yq�~���nǗq��k'�o]��}�bV�,�xɍ��t����J �0F�;�Vy�ʃU.���:eezyR?2��񱴢T�x�q��<K*�W��ՇW�ƞ7���H2��|��.����\S�J����g+@P�{@I�ǵ���a}�bʅ�#�X!z�����m9��\�1����w[н }�d!r`��@#���2#����9�.�ikW��{)�=;�C,$0�,ì�f��РP,ܷ�{N��6��h-MB�`j�T�a}�ȢR��65J��[���l�@ҏp����;P����	D�UT��������ک�$�@U`���5ԅ�Fa�T2���#C��^��z��lgҖ)ip�o�o\�������אS�#���G�=`idA~i>���^<��Atm����E��
"@�BαX���p|�&����{3
s�`�����x�͓V|��b��d��� ����<�.�ö�4��Q7J�D-�:�l��u*/��	�m^0�S��Ղ7a�)��Hn�P$..�aAFyq��()+�E�=��/�u��_��J��ȶ.AJ�U�X�@�W*�x�X�݁��=�ځ�̆=\����0�l�������?s��x� �٣��]��`Hv��'R�&U���2�-6���U���������¯�(��G��vLf�� %!�V�ߣǶ�hKi�8�.	=���?q�1�dB[�k�1��nqz�t��f�ȃ�q:�p�g�I%�%�"��rԉ��~F��t����$C(�Y�TUe5�lS2<+�
G�E���7_�o�!�*�S)�*��콸商�t�D��.AUq(���u_�o�!�*}��GE;����y���3C([��sS��B�--���*z
uCV�W��pcXcO��n�.�gq��k܇�V�ھ'#
Tޅ��!7�T��ic�+�`�������r���\֪`�f��g[�����������8Z��!ՓCCB��S.� !;X�򜢝 \Cf�Py�P�Z��~^U',�����q r�����?VL�n�Y�f��o������E���}�(���6`���x|�㸤�%xh�C�.��u��|�.�$�����n�u�p����>w`I��h�SFL������g�Ω�����-�A"�X۴��$WĐ:O��!�icj�s꘩��m�X^�'}?	][t�2�Z�⮉�ﳫ~Q6���h�wy����Q]��]���o���"�;2v������X�nQ��13�#2�K��!x�(; ��
�O�sp�Ew�qpc�M^�~m���`ƚj��0�#�cHP���k����8q�з]_��"��{����R��i7Pi���I���9�o|��Z��M[�2����%|�G����S�#�o�0,�q0fl��7�zW��+RVH����ݯ����'޿n��T���á���Nd�����`���/��i��@켴��2�Ir�֮xH�7����'�B�
�����e��~L�1�Q|]�����:��9vK��=��Q����>-h�ִ� ��2|��K�e�_���v0��(DGDc�wE[�%��U���?��-��:{>a��a����x %�Ѩ��O�;�ޑi���Gs��`�AaBVr�ѵ2�r�<}~�Uu��a*b�Ǌd�|2Yps�����3YEY(�(�]�܅�t�wVͰ=ǚ�w���;��l#\��7pѾ�Ȧ�Z��P��`~I�q.�z]؝����L]۟��F\�ٟIկ��II�� c6 3�݉�r�T�)�*<Uc�L|fv�T
c�!�����d(T�+Ġ��eg�|r���B�^�]Ǳ���t�3i3\v�(Ԙ���Nݾ����y;aG�>���QC���g��?���}%��m�!�*���	6�y�%��#-}���ޟyڏh��2��)��9������5�Cn��p���Q��6�'��Uٽz���w2�����#Xȉ�8x� �E�CǦ��W�.�߰�STޠ�Iþ0�C݌�#�:�v�Y�> ��+�|O�{��SŧХy�%���#��֍[�.~ʚ)���A�JH�c�����8�X���T*P�H�&*����t5W�D�|�x���T%��T��G���8D{��"(0���_�!�-����1�����v�ҩ-�C7�J{e?�#34���%�����:����Ɨjx^�������@���F��0��yhmm��8���*-Ui�JW���;*��Qi�J_�t�J���J7�D&ĩ�^�?���:��9'գO�Ŀ��K��=[���}���£0�������eʢG����0�82����R!"_�b�{�\{+�-�cP�A2�M^9/�x	N�hL����n�!�(=�hU�Y BU
�a�����3�}0��F*�s]�J�L�0���z|���Wt/�6�5Q���%�0G����G�c����o�wP�X�K�OR�De�={��?#�(�w�\*q0� >��1�������?y�H�&���?ŧe��gyO�Y�T=��JGM�=*q*S��I3�N������*�Y|�)l�J�28Ց<#��c=Ztx�@��~�@����X�����Ú�ܨR�蔳�CMa,�fA�����J����O��ދ��#vO,ʬe�zeW���iX�jQuq��be�V'�`�XYD�iZ/�De�d_�i�@�Tl�B�7�/޿�}Q�OY=���a/�����O�(�Az(�3jYC(!�w���{�p���
ԟ�{��A#f���wQUY��K�?�za�8Pt �W���jEA�7|��t�Tϼ;k7n��6R�O]bB�b�b���D�Q0����i� ��rw<S�%0����.Uq�1UЩ9�R�]'�R���Z-�y2�/�o�Ȉ�*ǖ�6r6.TK���P��1ߓCݗ����]cTcs�B�H�y���d�:�����l[�ou�5&Z���Ģ���"���35V�*�(ű^*�R�^H�]����^л.���r�~�7|G)!}�R}E�*��	�n�z�:��ϴ�|h><{#�[�Y����L�H�SůD�V[e&!2��F=�rS�Q���CZ��B%�l��T_D�U3��S+�_�����3�\����9]R�]�ꋨ�LP��'�����!ZU�MW��v��U������>�X�e5{�@�������r���(;G��uV�QRлRu-�bhѨB!�ԯ/#�S�b/;;�O�?IN����1����hJ��`��:{��P��%��H�Q�e��G4GV^"�#0�l4�!��ZJ�aؖ�3�f�]t;DDF���G����8mvR���=�*�Yh3qE �@�k�%�^�S'�`�
�i�\�Ż�|-���Ք���O��u^[eTWB66MC�bٝ�����b�WS��,���ƾ��[.!cƌA��.�����ٳ�l���F(�[�RV�/��T�^sFt��a-����7~���q\z|���-�ubF)��J��rF����cD9~"l��D�xB���p%���އ��t�L߉��]�ʏ����>��c��	ТE�/�b�R� ��e�5%��չP,ڳH����k�]+=�Fٴ��ݪ7�Zo�#�3��4���$H���������R�	��TE3<�#����q8�u
�6ď�G��8̭���-[�g� A���+��|Q�J��w�)*�¬�+T��ǆ<�����o�|#�Ă�1r���&<��m)Mw���oEzDU/����RQ=�T�Q�Fؖ���6�2s�5�x��q�]w�];_;�{&��?�ĵ�u=����H=l�X���e8y��jT{02)�(b��6L3�I�y#7m��B<d=�S{T[pӻ�0&�1��7o@�f������M/L��}�Q����LW3f���"NQ���O�ʈ)����%L!�ڝ;%�?��O]����9ZQ��'ܔ��.��+@Eg:�,w*�h�8T�5�aE�u�!�TG�B�B�i����r�G�����(//GQ���!qʺQ%-�Ҩ���E����4�A�����@:�?��S����S1�#�&�,����12'�Z#ʑ)�A8hb�#�������*���@iY��ć-�՚��eŒ�7q݈RI���2*-/�,dJS9䫃x�;��0B����:�"ʱ�.0�e��%��O*T�f�U�ꓴ�Kb}l����L�76:��.��E��P[�n&!.�1*i���G��sLut�!�L�H��Ӗ�Ȝ�T�/�r�J���>�*}������œ��fH����G\�Y�������!1��9�O'q�AL=~]�S<�y��ߠ��S�m*i���G�:?"�1���D�^��]s��@<�7Fu �����]���Bz��SU}OY���<ɧb�/!��h��<�y�(G�Mh@�n�u���:X*\����!�P�z'}|c��!-޹7�sD9����~���-0�C���"�"E��[��B�$׬Q3�U�t�i	�ԲuK�N�:���@4o�AAA(++Cvv6���*���|���}�Ij�?M��:[s�|�s8�͢}�0l�k�(GȀk�s�:#���J5k����ƞ�=hפ�\�$F_0�{�$m{�v̩��w�yUUhڴ)�|�Ma��/�������᭷�³�>��C���a���9s&���sG�F��~�K��/����ywi�En-����$���Q�:ܢ=�pWpQ��+O#�Sq��F�2�d��[#o��k����lq��j%dʾ��3g������K/���a�����S�F��4ddf`劕�	��%��I섷���`I='vء�X�D�}3A��
�P����	G\���le��Н��/aҲIHNOhsҥ�DE����ަ8�}��܇5+�����;�Y���?��`rrs`�:����ailxPq!�~��&�ԩ,�Z�?�iEQ��5��6���b�<Kkl���k�5�*S�~/��!�޸ikW�xCYy7א*T��9�g\��"�޻Z���7Nǚ�k�(��X�����!wa.nn{3�_���㉿<��;��|)Z^���]�՝V#Ϛ'hm���J7��F%JMcU���*�Q�Dg���vl<g��g�ʦ������7{��#����5�{��H:�d�/n�+�ܴ���r��Y]�;�R�N:	sw���V-Z!�$���Wv�RB���6�^�(�7Adx$��t��Q��Ъe+�.���2E���d	�5�
��"�bS��J&�<��#��mC����As��:�"vDk0����]�NM;aq�b�p��ӄ!�b�!�x��J���ܔE(��^�N�I:�ܦ�8�7e 屨V!gf	 �?��'+�����6�-�kyߔUSЪq+����%�.���=_9�8�G��ͻ7x� �d��aWꡨ�(�g�J��8U�p�|�q���[��)a� ��Nv�������it���٦NG���!�Y��Ғ9�Q�t�Hq~��ĉ|;����*ˑ�gXN�i3l3PQ`��u��fi�m�l,i�ò?RIo.���윚�{�#�p?o�>U��ŧ1}���kjZܔ���9�}Y-ڴ1d"�Ri�Ƶ�[��D��<�z�1���`���56�����m�lf��BMm��_]��$�6�S������L�N�^�>���g���:!���Ϩ�!~F�3j`��QC���^���>i����He�$��]�������S{A{^:�8ӣ�/������}���5��ξ/�l�*I���)�Ɛ����z�=C���Ʉ;v�V�B��7t��E�C��w)�I�;jC�O��}���N���KE)G�
Z�gec��3�Z�BIe	�S�e7�Lѝ�-��;���_��*g��k�F���t|���۴U~��Sb/m�HB1mMߊ�]Ǌ�����F�S�?�=_U���Sj����(r��z�{/�;N�xS~7S�zn���-���������J��QuS���Z����S@E��̝��	�s����BD��
�0{�lt���� L�YdGtM ����F�cK[rKr��:�%�/*/���G��v���U�g:Y|R:Uz~:�=�-ڴh#ռ��}L8QbhId$Z�Ӳ֛[
;?�)^�<��yV�ɪ!�m��)WO��~���V=��Q۲Rsˑ�8��=��8R0�{����͒�Σ�^����3�ߞ���?}���"
USO��e�T����M�䦭]�#*<����J�шc/��v}&��Q�Ne_����ت���&��?�t�!�!�~��N9���18z�L]��������v@ǜ=FH�O��<͍A?ɜj�,�!*iK<�Ŷ������=��0jp&⿦��&�����x�?3q{��epD��9Wb2><�aq�`��˸�Oy�����t~gK5^ӈ���qz��!��&h;@\�3�3�ս�[�3�ՃV'^u}"��҃��zi�@t����kCٙ	v�!�Ws��xx��������p��0ޘ�a龥���j�K;\*#������S�#�	m	�X����)��}9����B�6�5(a� v�>�����Ȑp� �9����Bm��z:_��)ʞ�y��b鞥�gS�}qŋ5��?���ؙy�D؎D�=���ߩ����!m�cO�)��v�y��Җދ�Gs�����A��g��?���50���;C�di8�����8�rz�f��`�U���_v$�WejUq%�C؎g�	0�w�T�Q]���@�B*Q�Cs��A��������Kv��?��$,��˴8�G:���8Z�c����>wFs��n���Î\����X�h��du3FAO}B�V�=^_��X��<�e�����%���A��&��w�#�ic�����W׼Zm\g��ua=υ�9UG� �RP[���z���v9S�������/�x��	o���W��_Y�
��>V�2���~�+�mG�-=���q� �;:
��X�ܽw��uG�a牝��E5o�<Q���]1-a�xUQEMm0�]��w�[W��-{`����T}£2hẄDu&���P��(q������q8Fw-���죢�	�#��响�kw6O����C�����#�'f����b�>��9�w�{�?u\*������ғ�G��A�kk_C^a�0IN��~��9J�Ν;��\Ϟ=ŧ1   ����sӦMزe**��w��&`p��=�ҽ���e�H�K�����3�Z��x���N�o��%lY�y%��B\��:^reHp-OjZ���fq>��8�{������"�����P$.�Px���C����5��9N��"##q�}�aĈ��n:*�ջwo�;�����㏱}�v��L�S�2���&����b�ƈO�X�ی���xu��v���.��"R����� i^��8�r�ɗ�^" ������#;��ud��U2"��|���B>��bbb���ϣS�N��[R�{2J*c@Κ5.�xߊ�+d
��ȏ�q��_{-�2�0q�D�
�K{��?�E^A��\lZ��;�pb�^u�`Z���繏�c�ک�i�@k�}t`ai�$a�A-=�������^E�Y���TőAf�)����	��GyyyyX�z��M�y
���oFee�t"�o�C��ʊJ9���W(Lӽ����#��!|8/_#�b�`��� ��A��?������=�,ggS�؂GO��A,��?r��99+���)2F��q�{�GFF]���S�������G�L��$��Y���D$O�~N�˓�x�έɶb\��o5vY\7(��i�w���?��#��5l@-����v:|�p	Dp�ą�u��=z4>��3�7��<��l3N]ta��6}��-����"���CDD��{�t4p�@�9[�w֩�-�E���`gB�����$�GA�y<���&�gCd&7���M�_PNN�������2��?��M0d�޽�X��#�����w�o�M0d�ΝHMME���C<א�+}��,�3C�}5<9�h�^�R�d<�H�C�T3�|<��32���ߨQ#$$$`�ƍ8g��i����x�(GE�a�Dr� �H$�RR��7�q@��F����y�I�&���Lh:z��~@�n�p��7��S�P8t�й�ϥ1��0���ư,���f�������=u��v=��A�����L_3]�@�I%�ݿ����0��ɂ�XCD�0o��s6Q~���8�z���T�8��Ĩv\7�X�6m�D�sK���(����gGM�Ύ̀p�n��Q���0���s�Fb�-j�o6?�He!��;4��6��"��߸�q2�h%��zh�}���O>�[�n����ѧO�0�K`=���=�9��o�{�(yFz��F�y>���@�,ø^�'������B`�������d4�k�k�?�z:����e�$�"@E+� frԑ.�fD`c�5�mq�΋���$9::]�t�MGEnn��!d�W�J=۸��$��̟f�T{�W��+_���K1.v� s�k�B�/13���O�ag����v��ƽF����Sa����y��������m��1���i%�x��뢻�8�1�K}JI/�^�ĉ�ϔpSϛ�l���������Zyh%n��A>I�� N���'�_��%c1Λ�čZޕ!M�@����HaX�a����dAt�h��O��a��uoH/��at
%�0�|ߌN�����[�Q19�I0�K�e��?O�)2��ȅQ"*,Jv6^�t�w��Q��ik�刅�S����0��Mq����<�5{n�sRY9i��CX�{�h�3�̚3l���_Uv���A���gb(\��^�)3��!Ft�c���g�5�mD���9�����:E�#"H��h�g��9q��K��FǿR��K5��f�{	�K:G|��d�a��,?��C�8�?�6QPQk�sj���y���O~�^e+�j�gJYtO�SD9���������5�u-�~��21-����ddV����;�p&�Djp&��v/�QB���਩sdk�7r~l~����">�@8NA���V��#�w�����v� ���@��x��3�'��#qD�a6�    IEND�B`�PK   [x�X��"�IY eY /   images/42bd9711-1b72-4047-a3d8-ad461b8cf403.png��e\�-��{p[ ��[ �\	������%��,w����^������ef��7�5]]uΩ�0%i4d"d  �&+#� @�  �lD���������@��!  �J��0<1@� јUw���� �~��A�,炳�W9���O䧂;>���o�~������*�j5#O��y��Zm���|)�i��;��׷�9>�^r����y?������|�
\=����d��ִ�ԇ��Ȍ�l Ix~���6�(``i��@��e�4b�-��\�N��wBS����"D�^���_ku�a�H�c��ΟK�_�wYC�Ѻp���8��& I���5�aǵ{�޴���b��l�/����䍚Ԋ��ޒ�aÖ�¨�w��Ce�R���r�AüE�Wq�������D�L�����mImkI���w����c�}m��à��r��?�;�{~��IRB�'uϔ��4�7��M��+G箷d^&Y;����_&C�'�Vk�4�f��o[q�(E�����5j#��a���ލoI�����jȓJ�	W���k���$F��v�մ���5R魍�˝�\�M�N��VK��+�>��18���Uw�۵�d�f�O�_���<.��k˭G��9�[���w�U�4�ԲM�py��A}�U
?xP��rP�(;p�-J#��銖 �ixLD#=A3~�|C4���j�*!Ǆ#��y���7��v�K�#��G��\���� �4���B�8�A,����R��@�	�<Sj���qW�|���)6��
G�fW�&gL���-/��-M�D4���"�(��@�u�hD#B,�2��F~�-Mo��×}j���n�e��F�
9�y��rPL�"@�*4vO����1�̲)��;9v<��s%�M�|�.�.f�*b��j3���al͋�58�Խh���L.���*�����Q9�S������-�l�t���D��6���.�A,6�����z�_X >j!B��!�Vxܛ�&A��V�ˋ�*V��~U��G��1q��9l�Q�"6.��Xg��_��;�6Ԛ|Jȉ��m�ұ��;�N^?<n�>��&sb���-�����������Iչ?S�=]�V�y�w6�ԍ��(e�d���`��6^%Wo(�]���k�V�E�����E����ңm?��-û#\ٸ �>�}�����q�����/}WxA>ҏQ�~���$9v7��4����D�h{{P�%v�ۿ������o�-k�_�8����<f�h����̶�(}܁ ��$-��#�S/�.w\�way��O�^��Bl���[O=N]��c��?��H�`GͿ�����d�b_m����J3�V�_����1O�%���O��:]>kj����)��	6� 9��h�~�,�~���Խ�q��|m�̙='�T?�-"����dV�-��M�G��,�'�8׊<
-����^�%�	<�V����J��׿�gO������������/r��[U����8�$�cLf{�兒���_$]G@�H:�Gm5\ݜ���
�&*9Ǿݟ��r6�rKu�TNڤ�>�%����jA�\:�������R��Ф�|F��ᝥtx�G0fAo 8�M�����僰_�F��s_�b�Q.�'X-��
������/����E&�,�;��ʀ|����S�ѹٗm��&�I��d�kE{ι%�����*S�|��: �a��O@I�s�s��Sҵv�j��b����O縉�s�\�z���C[�%׊���kL�����������|�%����B��O���d���˰d4�:���⢎R�e�������.�[A"���e��?
��
L��Z�?�{8�����l��%��R<e-�Bu�0���z`~�]b^�E�����vhE��{9�m��y�nϩ%�-���N��y�}C���&�T��ӍBw�*��ȇ�`2�6&H�+Z� y�á����y�"^��e_z����s*k͖��U�5����G'4�NP���L�;�����<֯o������q��W�"Գ�l`O`�G��q�b.����9b�K�zx�]��r��a�V��}Z�z�Զ�ZC_$����f6n�GZa:�9jQ�	�$[�GE}��[�������� f��MRӃ_c?��y`�C� ���/�3�2eg'�Z^���mob�xH��E�WD��3Y��y'�l$1�Z�h�m�4F3G��RQ���OO��u���Y��n/Pl��A�X_H�]�m�����>��?��/@����Z-3P�%�̯uRk�T�H�����P8y`���Ca�[�ZP^~TJ궴�Ǥ}aY��D<o�H���t�nr#1�Q���'�q FRۍ���QX}.>'�g��R��h�)�-^�739��'6_M��
����tjez��`ԡQc 
H)Ň`�k�<�� a��On�D�,������o�^܊8�㈃�#��b��a�k@cї����S������]ZQ�qYڬ�h�u��|�}�~�@[��}iފ,���V�q<�D9L�B�y��D`�#:j�͊�@0���m�ș�.��K�����z1���� z�m��n�b��\�� !_P���aM�)6�!X�pJ�.����{��3n���/ʲE�J�Y��W�_�L�d�h��,O����=��@E��2��h�2{��AקL��V��bf�Z�?��Y�����\�;;J�lw�\�<\ќ�L�+z���0 َ��)��$�S?�n`��lW��m��M���@�g�����f��o;J�6��������5X��뻈���t{�v�p�B��Ll��+7lkD�\O.E?�6��|�a5�dZK������]��@}���EI��/�9qk��N@o�Y$
es��I�+F�����U4K��-	��c�w���~�X�����cM��:��ή
v^>�j"��<�Y:�������l��5,cf-`b��ǭԯk����)ÎM�dZ�F*-{�X@ɹ�Vju�Gg��"˓DU��W�0����k���Y���.������Be�����?:T�O�VI���OOO��������U��.�W�q//
�uu��WTD�t�S�	�����|�eH�s-����/�4��ٽ�V�y����6��c����e�&qt]���xy�%yZN����S��`ՙRC�O�ޟ�ó�C�3���ܾ�Z�Vepۢ�q�"��<RYnUt�ν�v7��u�x.����m�Ε����W;�Ț\���%L�����몫I��z�"�ك�77��(F04p}��Z���}?�ՖX�d��mɉ�*�:�����*�:leאs	�up�5����R��/q��WZ�&��^�\SYUQ!S�h۩SRe=�ۣ�޿���Ȱg��Fۻ�~���l����T��.�5���̧M�v�msZc���7ww�G�Xb�J�r�G��IwK��l �Ӯ�3��('c��F�Q<��(^�ۣ��y��Fk�U�۔�jy�� �X�^��xb���h��"�|������b���9�s����n�fT~yu�U)��5�?(�\}�����RÞo�#m\T����c2�ƟN]ݱC�	��Y7������y������� �
S��RL0
TL!>��6�ɱ�0w�J@l3�in�u>U�4	�A"rwʗ�	�P���ԙ-d��T��/��$|��	��k_>0����_��'�u�'�ؐaZ
Y�ۧ{�3�f��O�M,�k�����8??��Uk����~�gd<z�,E�:�Z������~kV�����%�k�>[��F���¶09JS�@��&W��A����x�2��=z���8�*��8<�Z����7�C��J��%oE0$v!?N�܆���"DtxVw�t��V\�~�z�׿u�����+6|��=Zq��P^\K����>30Q
��F��ۭ��7�I���da-:VG��e-�˒�kv��,��B���}	<�'m�`������)�땏�y^}�:�i�>��?���Z���w�'��#�T7��tT.'�m�O�i������~�Ͽ���ۧ�~ ��2���b �E4��?ؤ���[$�>��#|�d C�w��P K�$��*�s��7�	�._�®��:�0Q�8ax����D�j�*T������!�Ժ��������6�]EE{W���mH��Q 8��F;!�V
�dv�?U��T(�����z���:��3B�d�G5�==I���7j��zK����/�p[��uJj�z��^��d��XdRe�m���J@��a$�7b.�ϑ�!��%/W`Nd��B~]Vշȹp `�����~�`"���)�_O���MF肠�,k�h�a��x`������N�"�+�bΩ
pQ�KR<բ�<��o/��SF���J�X��4-ɍ[�{��A�]?V�0���H����i�4��|����)pY��Q�"703~��\>�/�\NI`d=oa�-OO�F8��t��D�9�<�'S��܆��8y��=�=f�#hy�|M�뮁��k���R�VL7���`lM���}2��!=�n�?��ΜH�繁���2uf�o����$��/eJ�n�!z,v�G0nok� $�ew�c�5#���ikˉ���Ŵ-3I�ihR�h릢Q���%�3`"�B�DD[������a�|T�%r������+W��Wօc@�����8z�N�G��G�**ܡ��.�'��-ϛ�(���d���
�Oo�0�����k��+��8*��e4��nZ	r��a-�T��������{?��z�o�a!��sB`+�|�Z�pů��r�1(*�2n���N�}�W������_�R�q,V���,�R���ItzȠ���]��0Y�*S���hBw�/��|�*sn����y�C����B:�Ym.Ϣ��o�!
MLA鉨�CՆ�L�� X��pۚ �F`�w��06������_�Z:FI�Y謨v�_Y�c��n1��ϡб}b�GĴQ[��~����^���)S����|��/:������q]:� 7*eFD���������<�r
�����v��u[=]hu>X�]i��[���R�q�z�C�����l�����J�<v9��h���@��q��r:���'0mN��ʯq���أL�K��Y)09&G��wd��8�Uw늳0��!bC����)BT+|��u);[�j��1`� ��&tNW�I��62΀��@WEV܈'�d:�b�xּS�$`y�������B�QBj���J�Ť�T�Ч>A}��Ak��>����7,,h£CIg��	���³_��R�06���"�WO�"Ʉ' �$A}��	���\�p��[o	deeƫ�<	W`���##FDM����C���ȏ������wS��s}��Y���z�7��i6g&AYd�	l;�����S)���_��2Ca@��O�Y?���ɸ��ƫ��r��+�)�|��m�~��JG���Ƴ#8�c�{F��h�rܯ��c8�#�k挒�t��$0b\�@�v�����8
.݃�Xwā$��ǋϵ�3�.�L�3�|���]\h���C�(9@�N��n��q��X=d��&�;:��F�V1��u��,��rB�/1�t߾wm����U�(�}��$-坴�jw�pk�Q�J��jl�o��Viяk��$Fxm�M�]�H������r�}Y��oP�G���
��iEjof��'U���[����6¤
ڻ/ (.���W�0X��x����4�	$�IH0��o:Deკ�t��u��%�o+�ԣf��d�(���X+�ˤ��~�<�n�q$?���|��(��^s����Ӳ^�}��o�=��^5v>A�t���F� ���EC� R	���+SZ�"��+�_H�%͢g�@Y�����G�:5�g9�:���k@k��G�:K��.檡��'p���(�pj38辕��J��o�+������������>8�: ���n��=��<�O]�L��}��i0��`~��7���؞�/����چxp�?Zਔ:���� ih+��0I��R@��5K������yɪ]{�3<�f�:KN-s�U������5�r�P���'��ŸhK�i�x�ҹd�>���U�R�g�1�qۦ�i���s����P=�e���c�V�kO�읤FU�w�@�Cڂ�;���!��> ��P��'�"��I�@�<3�JyJ�Q0e!�3��$HD�$L�� ����Y�����(a1���;�Yn�&�A<��^?��]ݦ��,��L=�5�|9ЂOS�#L~АQ%��~-d������C��5F80�`���a끏��핎�W �R�v;��n�^EN�s���Z�����l"L9�9 �,��cWrw]�yk��i���27/��{�H�s�ְ��8_��
1�?+>�Xu����A{s\<��m�|RJShQ2����<ؾ4���
�7A�
���Q���A�YX�P5��Q8���/@Ze___Q&Ǿ��R�C^���RU}�]I�o~ïUC8�p[��"��Rə��N��;8І�郋�,��Sռ{�,��^_D-��$�FU��2�>�����UQ$x�]@�Դ��V��v��bU��#O2�o�����?�j���Q�.$C��l�u��c��7e�|�9�:ϯK���S���AY��
a ȧ�k�Q,c���^�_6��D�����D�f���UPqX`!��1��!jF��yd�T�>�������l1�xy~�~�ە��.�."!��A�ޮ�5�pG�ؒc�7&<��1v���#�4˳�����~_��!��������U@��yT���c��K��,�s� �|�0�{���ֺ���~B?[ȬiS��cҾ��{���� ���75#Ŕ�Ւ�h��HOq8ڴ�Y���5�5?A��xS+�5�1��<���9�O�gW����r]'E#x���c͡a֨����Y��E$�;L��e����eꙛ|��L�p�/���F�Ij��ڝY����d���(>ٖ�����(���3�?C��?cr�2p��H�m.v_���7�y.[w�����˺���gw4�u��������W�a�Tq~�`���y�%�0��	l��5d�����Ǆv�/�f+,�>vf�i�BW�!�Φ��V����@pK����a����P���(�h�c��,��A�L�)�mε��<nKU��>��訍�(�3�=Dp��Z�F����z>K��0�Ц��L ��Q���-WCug�B�y ��rt��j�bmqh�#��U�h�*�oo7�������mΣ�G��qJ�u:�N��v�L2��	6{���il���:�t�?�c&LS�
#(���9�׮:R+�j� "푯��&s��2�O{#�}g
e�|�36^�ls��ը6&Xk��"[��Ğ�]@��C_(��M!#l���L:N:��I�զv+��9sSMwޮJ>�k@�"4nE����]���4�f�Z�&og~����;��!J�W�خ�|��[��@ ����+F�����nJ��`�<�a�rm�3 ��J�ޮ��>J
��)$y�a�ǩ�s����ؤѭ_�Y׼ţ��b����S�VMlU��ʲֳ#Y��|�$�d�n��bj>�VS��K� #�?����%N��+�����)V+$�R�5������]�������,�W{������G�"��u~�����5��*񐲡���=b��j;N�:�#$	��֋�G��!!�9�Z�Y n�`ic$�r�܉��p�D���(������G|�6�KJI��edI�^A�4�|�i2������jI6��;���c4z�3>Q��+s�/��Q>�a]����T��FT��+$���F����&m�1�U���ٯ^g����Tc0s.�۹[���X���}[̹�@=�/�^L�.�sW� q� ���6�2�P b�|�������`����{�j��2L����T1���c��ߞ"��n��}��,��Q�b����UC�A���z�H� ֊����me#��	����P�Χ��E���
��A��t6e\L��h��:h�Ԅ�P���N 	�$��#z(�m,X��ͤ��J����x>�
%���K1z�H����~`1����=�Kȼ?����?-r"��x���En���8'EG�Z�������{�K,�6����aƨ���3ڥ���6~�����T��rT1
s���l��6)��I�q,���*Ċ�WZ�$����~�T@�ڷTs���~�X�k+���`S4�kϚo #I;r�iV�~ޕa�����
FàG�c_\j��F�!�_�Wt�U�1��c�?����KZ��ᴦ�u�p�9�r�f}/��d�3�$����J%����e�+��?tE��V膇����x�a �@*ꈌ�R^C��ݖ���h�։u�����;��c
]5ARD@!��<����u��<Py�m�u�ά@,a�X9�7�������w�E�?��xf�\��1?��vX�P�V=�K�܍�kN���Ӄ0���L��.�1j"���lvJc˖�"�%X�>�~;3�f>��.�+��Q��5���u�h�ӷ���PL��g\F�L�e�Q#'}�界ru��X�jn�Tac=hw�o��g�Ii�
ì�L���ўK0�$@o�������X�#�K
����e���C�B�=�H�M�ύ~A���ym�b0o��*�i�(�K�1ӊ��������U�/~ͼ8�/�?ԓv��Rם�u���w!O��*ΝM��p��⭮�靔���?�Iq��N��\Mŧ������6�O��q�a������`�|��:��tVi@�+�HI �s�)�˘F�{2
$�lE��Q1�\\}�e[ۢsv�N�ug,��(�T��
�i�ޯ��Z8"���G�9�������m� ���-�g����llV>��U��E��x4����Aq37��D~P�پc��^��v�֦�\��u�`"�>�Ľ67�o	�j>��t�[0⃡�d����8'_F2���*o��B'��npX���eٝ���|b���l�7O����ҰY��3���e\����aԗ��<' �}�$>�9�Ͱ�����Ԍ��FDD.I���jo���B`�ˁ!|������^F/#`O��.f�LCwr��t�#�Ӄ���O���Yq�vK�crI��}���l�:���NEv6�,M�ǻ���*��fb}�0L����V�	^���yu�&���g�!����������$	��Ws��|�Q��|���p��[E�@X����?6�c��3����Z�������nO�/4w�$.�d��ג�p�9�⩛5�"�4apo�ఔ`�	4�cJm���?==�(��%R��ҾO���k� w$n{^�H��c�R}�Ȅy�9�5��j�UBs'/Čb�\-}��|���ً�*Ϛڱ�y
8�06��,;�EW���d�[�~�����.����b��^��b��{�;�X9���d;ޝ�V#�(���UxF�C�N�ǂH��ʵ�o����\���2+��ջj����|�닞¬Ь#�D6<��i����b�ϋ��e~fWsQ��K��\3KK�j��m�04�H�	���].U�v�m_��JK����b9#dPi��9CԴ�^_E��Q�ժ^���tdG�w�hp]��bs�lѦBU��)��>�C:��U�;Ξ�YWw���گC�phёO�ˋ�~�(+O"���誫�|�!�+�p��y�GyT��/����^u�l���l8��Q�˓������{�C��\$�M����`,3l���	��Ήv�엻m��P��KE��*�h�*���`�����(j��)(�kK��kMc�-�<�_�c����F�e�-�;�E��N��Hٷ�#K./����7�����!g� T豟��]�4���m.���%������֐}/���=��*Y~q�<�Xu���gE�Bu���(C���Y+!o��������sSz���+��a��ٲx;,�@3G�r��^{\u7��n�4��""X����V�pd3Ič�!r0p�+S�綘�<'w�7/RP�St#9(^XX�8�7��b��k��naZ���^�ZKa�
�hhEA����'����J��`pB;�B�\FY@�����翄c��s�۔ظ�p1����Y�&�o]\��h�6K_�S&ĸ����Þ�� �xqE��z���l>mҵ��q����P�������+++�J��7��ө�j�}-,n4~k��N�m�d[cC���3>U����Ku�]����L ���h�\���jݾ��i�E�+�6�7�dH�=���#tJϽ4�yL,X�N��|�K0a�1)F��ql���M#Q�YhsԨbkC�F����t�W�l~�UM뺡�f������F���ea�m�Ŕ(�F�g�]�7F[q`(5%b�]0Ůu�C���At}��Ԅ�BмM `$���O,��R�n��)<��F�^��1BWC���'���v�Ĳ/�W[��~k�ʬ9�Ԯp��3e)-%�Uh">�]�!���|e�J/w�`��%��*��p���g>�j;�!%M)̄uh#3ޡT��1VF}�ko�@��-���w��w�$�d�|�xS۾Z�QJ�B2�0P_�`�U����g�Np�����7b��7��y]#���/�4wޭ%�(�_O6�rs�Fr�o�ttN|�%�f�קb-#_��r�����%.��r��Mg�~�G8��)�ܒR��V1��{cҤ$�\G��ߛt��رg����f��%R��*J�[�fY�i�`�A3ԤN�f�
k���N7�ߣ�@�]&�-�^ɮ����^�ֲO(/��	���"�%��y�:�6����C�v+��k�wȴ�3��iM�������b��S�*���*<�j��b��V[\\��-������#[k�o�$%�@�����;�Y���ş��N�Yd��/��l��@�@��ގ0N�>3̻@m�ņ!����]�֐9C����B�P�7��C)�+��&��p�l=�\��:B��p��/�|���[_l]{6��L�B�C����W���?0�eWz�\t��8�/]�eC�t$Y�cz�����D���7sUo��|��:�2��@2��������wל@�1'ܯ$lK�����4�$`ocߌ�!6�di����"�E,C��s����^�@�;�m=�~b9��3�w�i�)m�#3�Nu@�����u@N��V�KcO{��+�<��#|�p��ܱm�%�~�Q��.9ܑE{=ɽvq��4��ց�#�P�X����vaF�u8�����J;�Mk{YDȕ�{��P�JC���L SX0�P��`�����G\4.���A��U)7(�9c~Vy5�h�4�+�'��M9ZWz��Ԍ���A_�����*�6�a�$Jj�� ߘv��.�����`]�Ѐ<k�J�������V@v8��X�c9���`M'���A=��ں`BKH�e/`�d�]0k�����S�hZr���`�����R%ȁg���B��Tl�$n�������K�@�rߍ�n�Y�����ɶ0�LA�I~pe^�Bw�I�ZG'�'�0H0��:�N5�u�Jh	�Ĩ��5�c3���M��lL��=�[�MY`�����q���gDu��p�A1��:S��2�|"z�4ݦ���ɘ/��,�Ҩ4�%t���S�$�LO�Q>B3�NL��2_;U����=7֞������&/���i9U�a�x������"8�Foc�caEޠ�i�
X�a�v�x�]����O�5g~1�i�+�zk����FD��r�qD����p3���i^��N����� �����&�S��[n�S5�H�5ĒJ;+�"� ��g�����B��荋x�?��J�bC׋P�+�o�#c]!n"\
Kɚ�T�
�6�i�3��p�\}�פ�a���O��Ltg�D���-ͨ��w�,���2�W���P~j��$�N�vsu�PpN▹�PO-l(G�Ƿ��r��mQf�a�=]C��_$4&1�� �Dܨ�(qqѸ~�)��:0���E$��ZK�����|LL�}&@ս<?����+���?��A�|
Ke�):�O�c7_ ƹ�x;��4�� �BĞ�t��?���]M]�����/ bs��O8�����5�P���J��GnifY!���j!&"zr�&�5�<=�Ԃ�
�ISx������pa&�G������
uGG��	Zv�����ȳ�*�^��RB�Z�.�j�D��f�n	F!1�֝�3e���@VK�Dێ�Bl �@��^h�ց	��fw�bJ�4.��晌p����ٷr4jm�{��('�'�7���@��G°��Z��q+ip����%����Lm^� 1��ZDQO$"/���(΂��j�.d%@�aW���8��Y��v.��Kc�����>.�g�ܐ=�ְ�����&��5\k�
��}^�szB�9�P�UK��t4�s�����c8xg���RX̰�3X~���o�\[��ԶT�v����y�t�y��;�5�1b(G(�mB��K�7x�c/�X����ʎUP�++%l�|�NҨH8َ/Aǫ��~��e��H�,�A�׽�i�#J1�C$2�,$+�Q�@������T':V����$R�tZ����yђ,���Ԟԟ���|�c������'���F�{�wk���7�#�5 ���Gb3����i�DbwG��v_��~FI��TlߜA#�`ґ	��A�IҎ�3���O(��]'!p���g� "U�`1\�P��eu�	m�F�~�ʨ�;Z��vDG��B�޳"�ˀ ����E��4�_��U1�o~��65���{u�E��]�8�HD~��<�����oGycm�2�?9�!B�k����%6�,,h���8�?L�ZB9��ؽ�z�I����|0�j~��ށ:�TjR2ѽwR ��(��bր6�X��TD^;�Q S�V�i�V���~��l	�C�@�>~��Ȁ�қ�uDo:M��V��+�SKL��a��l�hQ9狅<��x�)8��d3�XXrhY�G���%��[֢�G�F���"�t�ON��)�S�5sX��db컗�������|��ɔ�����59�ސ�b�HJ�4�*Ej<���r��:���:��Vr�)F~i��q\u�F+��s�_�/�rN��U���K2'��2��������.�N�"���;��U�
%��T��v,�}�i&)n[�o7%��2A����r���#�P#���}h��4�%���'��P)��)p��@�Ts#�^8�st^��Z�����)�CE_u�J��E?�+cDTJc�QO4
�-����w��,T�2�;��R<���;W��/o����"�e��Ʉ?=t� '�SH:�O1��pjK��L��P�ۣ	eCI2�2��w�$�6â�T�H�cB��O�j���X�>���S����f0���sh���7���	��;���(5���?���/���3�ny��_σ,��4��
���׻eN)��3�6����n��ARw�����H�I�w� V?�4qJGI���SZ�T���������m�O�J����W{���<�+�<�C�?t�Z�AIA�3� 6�����PRb��C��j�W3� կ"a[}�lLKl75�'?��Y��u7w���;�}m��fy_��i�P��3AwH��/��Fw����18��C/zyX�u� � ��c�@���¼�E��ge_)�5���>�@ �a�%?��<��!�8	ikcc�Ņ�_Z�V*���:c��@�އ�4�A�D��%-!U`G	Zw���Y�I����8Y���3���p���!�,�T��獛�>�z�R��0��D���FN�����l>GJ�_��?�n
�kY
�5��|O-)~���!�7}C��HD��0��q1>��I�+�!�Yl����,���LMƭ��8�Bq�Lxb�L����]ꐕφ���|q��'��S{�c�P�׿�����EEu���8v�z�Ν�9�����Lς�_����ȝ7W(nC�z�����.�� �8l`
����yw�4�2k�P�NQQq,��
�����#-G����� �[�3���\�Ԋ�/2����c��gp�>�V����]@�
A�#A	�����^g�Y�-���F�Ʒ���GrlyC�!6���U_��`���Mafm:3��*o�܁����v��q8�����yVV35�}}��Wڢ]���S�����P�x0
r����~�ҍٔ���+� `K=�x�[p���Bz]�x�@�d�V �! �M�	��X���n͈i���A���E6�-�a"pH���cGB���1���L (�@
DS�.��t�Bt��5u������h�ll@z��;�h�����d�Z�_Ƅ��0�t��?ȁIWQ0�l�a�J���.�*�%���Hl0q���
�����!�Uua��S\��сDJ�����	?�&
a��t��n�No�y�<"$) �&��~	�.�ͧ:�	�f,�]�旇�Ů;�豶���z˸O�*���EG���?m����Pb���ƣz��<�� w=�BҒڀj��c#u{H�
��K��(Ky�)�6{(ߖl6dO1K(���d6f�|�>��r�e� ���B�}��4&��ڃ�4X[o1�w��g�.�A-�0Lh���<�*��4,"�y���'Ii1���-��蚶1�����F���]���I�W�]|E�0�{�dM��ᶡ6�������������~�$d0�����D8W"%b��[�R���3��|�ؽ�IM�6� Ɂ����aۼH�Ze�ؾ#.N�����f�@���r��s�
�hd(����Io�j<���zH֛�z@�ɩ����_�uE*�'�V�ap����h��;�~c�(���!�M)Oi�)gt�]Lxg��	���#��g�0��B��v@*f���0�,  �K���J{9J��p;��ì	�_�y#�@*���~�i]s4���Eh�����z���{��'��ݗ�����J �s�+�����$\sR���*���p������Y�0���d�,>��i����~�ڼ�'��=��0R��1�,��I`'�#f�`��CUj�S^���D�;M$4}���y�<��0�48����L���M�qb�����BJAQ[���a�4T�h@���e����Y嗄�J{��+�i9�%�ǢϺ_R>c�A�$ @�P0A�#�����s���vr6l�HPFP�i�2̸`�@�I:F�-J]-8�^�h�?a1�n�)�fX)
��5�y��UD�t��@< t��e�悙�/��n��i���@����������i��ԡl �?��BZ�mB���v�~xMDے�3|Є��;S���`���	�z>Ø��KK�ٲr�'Y�k�[`!t�ųK�P<��zK��:m㞛�0@���EMN?$����}�A(�V�����F��C�I"���BC{��$R��KQ�$�?��?�N|����xC=���ql���F�]f�tK������ֿE�9ת�Ϝ��T�i[Ռ�����|��٨gU��+��@ZV���Ģ֧�LN�fY��'�sSvmZ�q���Zҍ��!mx�w�!0���3�DGr�(d��(q[��,�ַ�Cd �2%�p�A���\5H���ZY1�l���Xڌ*t�*��;<��SH�j<�+o}���Mk�ە�1�N���xe�G%t�kk"�ՀSr��y�B�kίt�_$��oZ�T���2eG3X)~������84FL�k��o�-��wI5�d2��jB�g� j)����/"�kS�8	�UА�kbZ�K6D�ǏZu�H�\�hc�ɶ�8�p�}��G|)d�t*Ȝ�=q�'�yy�0��t��
�p��*�)A,�E!)�[�w@Bay^����$��we8V����B�\-� r��,!��>cH8M��o�)�*�4���8UJ���"����>���������`*��p��{�n�h]Fg��0T�3d�f[r�*"��.�r_���iF<�̼3����ƆN�p�������N9ݸ��ք�nI�2h����&~7�~�e)Q'�����{�Z�a.J}WʉB9���N�-��v��of��.�\���U6L�=�Y@�7�	杀�s�Uw6-ƽ%�4���@t���� �t���v`����A����h;X� '�,�B�E_���+iC�� Q֖-[�q"���f�w�}7�ꭈ���]zŒ�+
�3�Z0��c�m���)�!�2)jUs�>zu�˴j�f������B��*�'�d��� ���B�n"ɚE�=��ә�/]��c�/��b^#m��<4@Xw����X�,���*E���v¥tՁρ��'��`��e���[�lP�����h�޸� ��6@���qV�KX	j�����p"I����]��oo�9K�n���҇�p�g�r��C sbvG������h� k l�"�J��o����"���z�N1(��g?�g��فo�n钥�Ϙ1���-�Od�@��}�m�N��a�9�DGqgQ{��g8�/q�ೞ�Lt�=��eˠ����y9�H���̝;�Se"���{.� @C���+3���Id�Jh¢/sSv}����8��4��+���� �C�âYn�?��]���X"�$*"�� ��c��At�_;���* �&v*GG��L�P�&Gl�Xad���^����_� ��!C����f���������d`��X�^�#�Iރr {B���7�#m	�Z~�u���(�Ţ�@ =fi"���K����ԔT:� l��_�}���~�#,G@@���`1��*2��5��P _��H U�.p��1DO��'>A31�3v���B\_"���9܏�2��rHY��p9@��\記YAzB[@�]��tNY]��㡝���@��"3$ee�r�p%�D#�L�P�=��,G �����Ѹo���� ��� Z�'�p���>e���.��#���o��wQ?�I��aQ�,�A�(��K������Da�N!k.���������*΄k����Q%�����'��\O�>���4��;DlLD�C�d�PD�����
d���0�E�
Tc* �y#F=LM�^R��K�!t����ߩU^8�_���ԡ����ld;8��\>���%�\�!CX*�����}��%K���mRd�9��) 3�E|�S����v�1��M�N;���c��Vr�UU�q��X,�5���;bW�Ry�GÇ��XĦ��ZY�p��/D�\�n���|�v�,�3X���e¨�,�3�=H�'�fx�,���5D6�mao��F��xa�1�	x�&˜���%U%�@�8� g J����T ��~ɒ%�DnP�)h8�ԝC����TO�>��< � b +��#@�
"
�a!0���`�0��V}z �Tp>K�K�'��e|�녕��(���'��@���_�2;D���_���R�B�B�<����z4ˠn`�f��lS)��^ �x����\���� ə��y��S��0��<��nm#��`�g��r�,[�凫Yjǖ#`GHP.�.fݲ�	��N����-ā+�D��, ?p�a93��s�B$S�/�؆t� o\C4gd��k�Zok��40av�%�y�V�!�l�Lp���P�9��	���'�S�0D��Y��\���7�'(+�D��C&\N߶���YйY�i�$�Ơ��^��e�{Ǉ��$�Ph��b t��:t]]��t�eG�[��ާ�XE_q]$ٲ�g����6�+���>�H����O���d2"ݫ\&,˖/��"����&��>ș���(	Y����I��y�x%۱	pd�W��C�Ůz����f��ZZZ�U\�hغd�H��I����Y�P�*B[;��0�3AR�Ĩ� !��tS�o�ы!�x���YY'M Y�3*SOa��T����5ϰ�\�g%�@Xr�~�_�A���$��`��uG�����>g���*�L0d?�]7�0���`��o��rx��͡T:N;��T"�æt�#�Y���#��K��]�i�0�> [w��e|q�-9" ��p,�?(��^@%O��6���r��cP�h��%p
3v����I�Eڧ�ƀ	?���rn�AxX��R��јͫ|ȵ����8!vLX"$� F,�	�a��sNd97�w[�P¸zܱhi�����0�$�A���=���mu��5�\���!RF�@tJL+1E��/t8	���<W��\=��l2<8�l������C��R"�A5�1���7�ܴq+�{]��j +�D��^��v�A�|-&%S��{i�^�s?{�u�ԒR"%G��GV��Yl*� ��ñ��U.��LGw��;y���`�K"/q��;!�%�j� �=|���`-��6ᆭ�~��`�X1��fN��]�og\=c:� �taǨ n�Gc]L��ٌX:*�?��;CdU6C�u�P���U�r�0�10"#���zv�bօxqL)!Q@'�|"��s�� �@���A�lbׅ$Y�C��9���h��u��h�ȱԶ����p��jK�l+F�T�b1�J��uS]}Ŧ��9��Z�#5�x�J02���1���3�z/��+�T�!2c��U�F��p��X�N��	~H�S�9�1r� �����B$�,۶��dɒs*΄�un�d,�H&�,G�1T��e���,�+��l]W��eDp��	�ʻ[��u�2V,���2��v�J�V��<���s���:��О�1 #h^��Ndv%��ۯ,��)�) a���L0�%R�t����9��葿���珔L�����*��cQuM�z{6Pu�G��z���C(ѓ�_��z��)�Ĕ��L��uc2Dď�U�����aܕ�`�~�w�ل��	�$4ъe���
ڣ8NESFy:�	��H0a˲lii9�� �sЄe�\Ĭ�c�;N���=�~C��
��8.���d�:�fK0����G/`L�WʔN���!j�,��rv�֡i���Rs��<{�ˬ �UO���"4�B����5�j�אَA��ɁT���>���2S»�1�.��:���9��mS7]��[����J�]1�u��^&��&Ǎ�at�QG͢�.?���g<|���t٥Ki����%��5̂�b� <��S]����aѢ@�\E��6+��ܩ/�2(69^pI�7i���l�I�H��1:f	��94 �V�q�����2�z��{���%2�	x
��ߗ��) ,[���6)�(z��ש������ib�U�4ȕ�`�|���.��v:7Tv�Q���\�$SNc����k�ԇW����g¶��pH=Df͘�}�������"v����?�-]s�w�Pu�Jۈ��{��ldQr���I�g>�x�}�Ewu�袋��G}���*r=�c��k,J$�X��\YP��d�:���-s?F�%�q�m�䵰L�0a/�����#����I����t�@'f:��g�l9R��e�축M���qKȂeY�x�p!���B�uM&�u �6�_#��} ��ʕ�Qo'Bf����=�Q,�_i�r&#)����B��v�w�E����g����R���5�G�̚ <�H���{�5��X�%:`�T�x�G_��{tǏ~C�UM����2c̮���6-���L�5)�s�1�ŋ΢Q��y]��6:����Օ�ɠ:R^�#"��lJ�:��[p(��_1������:�LT�U�~�1��YO��@X>}�\,�N��H��8儹��>;�{ ���/^|vESY"w��0{��ݖ� ��;�@��]�{[0�� ��gJ������Jf�1И�V��#��Y@c���Y�0!�	�����~���e����2�DF��ش�t�Q�i���я?���wQ�WQڱ�@�Z9@��z=�϶�]<����(}���c��x<A���~�ӟ�A�=Y��p�CZt�-�y����g* (���
fFy (H�3�~ f����'�}�, ,�$�o1=#Ć��f�2��R��yB:���+V�8g���{��{ʐ�|#�e��[%�/�T�NF��Jv��F*��a
MES�Ҏ��Q �W����Lt$A��N^�������X�Ɯ��}�Di7����lJ���o��1C�l#�d$)Z�rV��fq��$UW5Q�!rU�s:}��̣����j��t���"��ck�{��0�V�����+G9�g�Ad������* ,�vp��������a�f��'�E$	;��q:���H�l��� �ͪ�m2��
�n����Tt�� ��	O&�°��̒�d�w	�ֽ���v�L�C�꥕+_���8Y`% 1�,8�����<��������_C���҅��4t�8:�������(ք���jiJ�{��;� �I���y����$�4�B�
��;m��! ���]�E� ��C��R2��H,ʻ��%ۈP:��6�Mv����7KLK|b��>�zM�x������;Fk�;�d���S�r������W^ynEA��7j_wkM�{��ә���+�k��#t�~� ���5�	��p�Au���/Ȏ�i<� c�x*�dv�:�7TQ�LJ_-���1�c�Ow��|�^x��`��SQ<��a�r�}@�1�2Ps�4��v��C��I���"� ��ҞK�!�b�h���`��b�����qd9�0�8���L����e�BLX|Stv[�g�.e�\	]�5
�lXo,�dS'�Ax��˖-;w��魃id7�l��zk��5)WtxBu�蚯1��M��5���ܱ�L�|�U��a�r�,���o��+�tI�h�.�a������������
u��N������c1*Ή{�巍~P�m�
��Kv/��f6��������X�gY1�OCԂ5)����Nd������M������0_t �2扦��]a����ئ�{���yf:�f��0a=�ד��L�	���g�BW�w |߲e��ms��Bn�	���N��BŰrl@��)4-�A�s�lp�Ż���� ����~4d���ӊ`�r^�����TXm�r��^87{:�w����6�p�	 �~���ֶ���@��ة�8]�gb`��5�6��$"˦X,B���c>��
̖#5�\_�,$G�kC a>L��$yn��qҰ���Vˢ���F�r�9+d��%s<��[����z��dG� ��,Y�+�rQ`�����I�2��\�U�aܷ|���*�[Zo�IuMB��D<E�U���dG���rF2L9��	�e��$UF�4�lBJ8$F�)�>�隱x�рa(�=�~���2U	kʌȈ���#�wf?�	���ʡd*NQ+ʫ9~ҴȴmjVG�M1\^��0_������`��{$���З,�o[#nu�Y�A��+�-^�'Y��%xj8�1(+���[�`Ov�0�o}�^la�Ul��>#	�		��|�6�%׍S�mQ$bR:��^�8���f�u��B�j^y��yWt7�I���ό��"�r= K��VObf�|��ÑL��,�@�� �x��">�qQV^�~������G��xG��>;g���)��m��.^����3g�L��/G|���M[Zo�%:&!cF��H-�`}M��{:9���C*K ��X�1x8�I<DT@e��ȳ�>�ɑ%яhf"����908�(�
�8O O@X���Y�Z7����]���R*N6�$�IɄK��"v��$�	"�!;
	1j&)ׯ���GG��<����;63ʹɧ���{aq�	 �^�&,;x� ��b�Z�[3�
�w7�zup�{�I�`��L�ӎ�d�d" $n��V��Ӧ��CS�΢�j��E�[�|v�T�([v�f���|���g�������I��?��o�C������f���M�G��yG ��4Y���Y:� l��T��)9,p���x�eݳd	�\Yn���͵i?w����1��������Q�|C:9��|"x�Rا	,�Ǳ�',T�	�׳a	`JN
+��4}��.��z0v6 ��� ����Z[_&�H��ɱH�5���SQr�AV���a6��4��5���;��wH�[by�Aٻ��e��LA��_�`c�`߷PފK	��[a�,�>�Uib� ���-XĤ
$�6* ̣M��/X��*�T
kO)j�4���jklNs���U�`󇣨y�Nd�H(�o��,Iؑeq��
 ��aGu� F=l3����^z)��u�]�dO�S�Dx������ ��^�L��^a
d�Cy�+�c/L�+;6k$ϳm��ŋ_0k֬u�i�E8�޺��LO�TrrG $�����9���7��-F	<��p]�Qd��4 I�![@w������h?�F\5�s` �k��H�P�����w�R0:���^��Y�G)J���ݽ�b1?�r�dU��[hŊ��֭.ّ*�.Ǔqf�G~�=a
��.��ϻ�`���X�B��̪ �U��g�@F(��} �K�g�jx	(@X��更����a�ʻXD�ʤ�S`�!>���Ѻ��ɶS4���>�S�}G�1� �xJQ]�pRf-��DK�UWײ��Na[���i�O~�LĂ�q�㫯��������9s氜�裏���!���?�C��ȓ�2������%��ʲ;������������>C���D~�hѢ���-grOo3a�0nn��It���M��x�Lx2���3B �� %F�5��7��'d��p�@�R��5���������>%Oh ��K"��@��������˒D�;�V��$iܞ�����s3E#u����􉏟O7C��%G�)4g�?�|�(���������Je�ʻ�T�	�re#�j�GH�~N8D++�`�>ɏK���m�4��0�a` @�[��6/ۊ���Nx������G"�륆Z�/�O��9��V�����^j�HS<aP4�@N��>S��z1��� ���G�!|o���1c��y���/2�A������П����7�̒����@`
��P�ꃄ�M�I$P�_�XX|Z�C� ���{�e�����"���-Z��� N��z/>L8��s �O��#�|�?|c�#��9�0ȊC p�]5*��[��Q놁q�:�(:묳x1��s��N6�mI�%+\p.v�����7�N�����:=����F�l�̙{�n���xo�^}i}�c��4���(�d�s��t���e�roO�L�����!�����E.����Y�pL�9����|W�����;����;��Z3��E�E���g>��O���sB�P�+_�_���DnE�]�x>�|ұd��J�ko��g�}�&�=�jFS*aR4VO�
R��sv�0������a	�����?�����3����d�©��������'^ G`ta`
�駟�~l
&,a�����*�u���E��p�������.���-J) �p�*
��˖�	E<"v-��1��<���]�7��Q�b�|������x���l�=�k.�M��\0�O<��xE/��B�
]u�Ulp_���������׼�y�vut��W�ڶ�@sN=�.��T��W^�Dg�u)�kMYu���r��� M����^-�(�����s�����Lh���\c _�/k �K��cy�r�+.3���}5�c8���� {����L��,l 8�;���;n%�레�K�z!���㑏����7�u��]���i��#(��)��D5{^�}*�YL��3 m���C��R�8�́�b��~.�
�|��\�8F�_    IDAT,��<��.B�d����?:�.A�����cG�O�m۾kѢE_�(O9w����kni��T��g1���/Pm]�|������Bb�͊sM �����(�P�d���=v^�f}�H�y晬A��/}�G(� c��C�\�&�r$װ��E�o:�����詧�JӦ��o|s�3~z�����ͣT���	?�
�W`���79����Qc������k�>��+K9V��a@v�eÅk��8�xa}1�3�%E��tr�i9@8��JU�-^|}��'RWw;-�j=���4z��w��4}�!�(Faf重b"�%�����u���>��>�Cd�������±���+H��ԧ�3H�
 �z����(�ɕ�<�(.�!�\lf��������g�毮����}ϙ?s��ͷEz�L�i~�F���g�m�z��'�̎�_q�nZ�P���#`D��3k�,�X 3�%�~�1��7�J��r
_���cP���Q�!1J�%�a3?8���*<iX�����+_Fo��53i�U���L�Wm���9�M 8J
��(F���~���AKB�B .��#����9����b��$1��Co)=����	0�Y��~��[(�襆FE�_�Y:�#�Gt��W�SO�Ұa{З._D�L��'�1���Xq���L;���J���z��N:�N:�L��K/�Dw�qmذ�/^̑7�x#/�8�/q��%��AV=��2�H_��@��������~0H��tJVṑ����._1��ɓ�Ʀy�#&ͻx������${�q�]e��	��=�^~�Ez��g	���� ¸A	'��1�'`(h7�
��2�
`��a��g�i����aA�q<>ñ-Z��� �qMLAp���>�������t啋�����A�^��&Mއ�{�u��GϦD2Fi7J�YEdD��9gp��q!���Ǿ�,  �曯����	�vwSuU�/9�N��<K����7��'��iͿ�2�c�=��7ͬ��N��㽝��C�����А�v/^������s��	'��}��?�}���e���׿��H��={�l:��=��;^� 	Y���υ܀������G�����M]��
Ѝؑ_/Z���Lx�s/�6r�[�ե�3"xISt�!G�	'|�{��f�2]dK�%��������L��w=='�PBBB "Hii�@��҂!�8���w����f�$� ���)�؝QQ�+�9m������OǓĐ'�u�u��������_�~����?DfI'Wp.L�����Z���p�҆��68���"|���P��r̄�6\�n����^��]{�n���q�����[�ՕU��R/��1��� L����,C}��%�9�t�}�*�rjk-k��߫/:5�y��g5��V�Ԫ[n�Co=��`�V��4�<M%��7��d�~����[�DE��6��;묳�S�����'�ֹ�q��8�Xm�|7������8�b�s-�n��N}���3�ל�r7o
�S�V+�T��;�ν���L�8���=fӚ�z:�F.: |��O�y�[?��g�a��s��7AB��:�!�r!�)��@]��Þ�|�K_
�{��;<��0e p^N'�fr8�c�%�s1~�bHV��ٮ�������Z��I����ڔϕ�nMY�w�r���%Ӥ �f�$O~G�?�����k[�e+���^j�&}����E���Ƥr��^zq�~�����7M��_?��_���l0fHS���A�!l��	����)G�ڈ#�y�����?�A0G��7q�y���d			"�t YH#�P���+w�h�r79`���4L��JWM�SO�}�]7�r�)�WE��o9j�����Ӽu�1�1�2�������^�Z*�IPI� ��TX;�� k5�5�����Yp�q@�^y��9���<,+戾��t�؎5��Љ1�=!$-�}�7YU�	�Sz�!l	�U���P�{�K��1�C��ɪTM)�	��4y�t5n���!~m��P��FᕫW�Ա�CMMe�}��5mƹJ���Jjn��[Kڴ9�|>�Lj��R�{�q���tD/%���1�Ad�=��}�X�17`�%�!�c��v�i�q���6��"�O�+����X�ҥ�}>8���Y�|ꩧ�y�ۄ��L���wr��Q��lZ����?��,"	^�a���ks�F}���U[#��W�X\p�/�a�e�sh �EP� :��dђt�+B�q�� 1��s���}��� �j�☳(�����\k���y��[3*��)��kX�H�������ھ����&>��*T�԰W	����vH�	0��s���@�ZHh̨V]u��z׻NR6[V:ԆH�\kTwgM�T����*�Jg*a�Ѱyp*�+~��<�i��aj�[�xm9A�7���G bS�N 68;�u�ĉ/���f�,0	��h�+�=�F�tWOwg2٧�y���0~Ӗ�����yՂ���I�#�Lވ��:u�8t����3*vcG��h,����߀'�^<������9��H?�&��q�{�F�5? 3�����/� ��a���X�`SvP��s�)�8kz��O�k���BO��P�2���k�(E�rج$N��K.�l��UO���x���P;C�/��C=��m�n7ftV�U��[�m�*U���ǝ�7��r� ���BoAz�I�,[�kD0�K���#����B�0���ի��;��N���I<'	Q����w`��8��`����ӟ�e���V�@��s�D�Z%c�s�����xío�i���|׉�d-I-��d���Stҩ'襥��r�������z��:i2:	���Fh/����C��6`�>���SO���]�Vs��	6c��m|7(�F��6M&�N���gU��:gRd�P!��>U�V�V�as�ƍW6C�r�@�Ƽ��kH�%+i���Tʥ�%ns�fʪVzTKBrjjl����Xe�#U-g��ܤ���`��ը�V�K�
[454(�ӼP 8�$���2�!V�����,=a�u�5��H����P�j,�v���k+v�&Rۃ�@���.����j�J)˯͙3gp����_^�pT�<�;ߝhmjU�3�7����2���5��g�5k��ES�ދ 錗f� "��I�-i��	=���3_(ڇf��@TT"`��k,���7�d ��q�۵t�":+��m-( )_`Ś��F���QBS���QGMP:�[����~!�PS�Z1�KOH�FU�Ez�N������6��Qo����ViPKK�����j���z�p>` ;��9	V�z��a��s��F[�3�ӎ�]̙�� v��6mڴ�z&��2�{�F6��ɢ�j���}Y�qސ�k�H���ܹs?4�E��ћ6,l��6)�I&��/Sa��u�X������MZ�|e�`�m:�"�N�0��d�j��x�t1�`r�Y�pZ{?h6�f�-溸� �����v����^\[��|O=�;Ö0�P*�6B�Wo��a[���
A���Pt�^����$`^�v�>���T쪅H���4jX�O�Jgq�Q$�Qg��B�:�ڢR� %;��)U*�@��G# ��w0�����vK�-���~�^"�LxhBÆ�]w��#��v];��@���8���xa���MM ��G[Q�"HP @�v���Lx�A���ͫ4to?���A����2h��*��:�Lw�[C��@��8:�Tm^���/t��? ��cE=���P%��% ��DG`~`9�&ta��"��7�!8�=x��xƌ5�(�R&�m���eU,oWKKB�JR�}~�>��g�eK�������Sg��!~���P�Q�+����ROU�nӬ+/�9�P�,�*�H�FU����u�R���������p?Ha_(>0Z�����?���%�)�6u�z�Hڊx^�s/g�b����Ŧ��z�OT��8�_	_m��QZ�M�6q�������	£6�Z�Z�91�N$�@��F1���+ۘљg���?!�V� 1�s99k�g9�ҀNq&�t �������\G�������;��@��a�$k��w0�2ib
z�ڵe�
e(�פ�/n��ݤ��ʵ�  L���(C�A��C���%�	c��֥�6��;ޫ����/D���`utI��P�I�r���l�`Xg�;|*.��5~3���RO|3���0��~z��:m��!8�� ��?f��W↹ ��~��6 �	��b� ��x�z�Q@�����Y�R�>��J�mI�=eU�5�(W�Ѱ�vM�0Qd�'L� G~��� a�t����g{@�(qu&�
"h�9;��N:�t���(�	;N8~}�a�U*t���򸎞p�N<����Vuu�fUQ^p�*�*ײ�
E|�N�g̑m7��=V5pI� �b��������'t睳t�{NUcSJ=���,ڬ<�k�t�jh�Z5�T�1D �{��f�@�d�x�3�Y5ϛ7/�%����e25�1U0�!|��<G? �|G�	��s8߬����^�S$������O?z��7 VΟ�H�Ά����	�E�a(��÷�'���cJ��@g)��vT#XG8�e1�D@�|�^�z�i�:���	�Q�o�p젣��|�>��U�nҥSߩ�o�'w,]�U�\t��y�8U��as�	1�}4Ǉn��K� �d�KZ��Q���WB��E�X�����O=�mۓ��#Җ��f%�ٰ�'�!2��'���C�U<d�3w�4���js]	���fe������������q�iq���^�Y���+l�؀c�2�5��+�L��a����$%��b���d��锺J��nKSk�xd�@�`��~m����(��L�^��pq�����ý\�Ӷ�s�m���r;8F�U��z���ߵj9�[>�����o~���8L�����qoђ%�4����;�r�A5���h��{A�%�s�9^5oH���r�r-|l�r���f�ϸ��@���������G��YW�_o}�۔���Ɔa�r�y
q�3�	c�c ���A�^ۡ�����&�l�^��`K���ڮ��u|/�
�����*��s eL|o_�K#ĵ���e��|�I�jI�M��娘��R��j�.0�t��i�5���BZ�YPt֬�5�^�g;��m֖|g��� 3���`Ψ	�^-���S�W�Я�S5������'u��oՒ�k4y�U*{A�-ﳚ:�
u�ذ�V�N���e�탩>t��Ua�'L�Rʫ����o��)S���C�S����>����;5~�DQ��'_P6S�=&���B&,)��e0����j�ؗ?���x�k 2��:'�6f��zTŰ��ͦN������Lc&<w�����>$klX�c�$!jDG�Sź�y�j-w6��^P���ef�d�8Y�%����~I�Ҡ]�j5d�}|��ziɯuđc�����z�����+4c�u���ܮD�[��2�2����U�wr(cn_�ܡ{�	$����+ֿ�+���pJK����Y���i��>��Y�>������}�k?Ѩ�o�-~��;A������j� L6m}g�N�c����v�κ��{�|?��jb��cL�ܸM�f���͛w��g�mX�������
q��Aة�����}9�x��������{�Ś�O��������#ںu�f�:O7�0]�����3oԶ��pk�'LL�)�4~JgJa�!ޗow���^{��Y�A}D=]���V�w�O�M?O�B�~������K�])}�c���'ջ�H�B9��-��Y�9
�p�R�o� ��c9D�^��b��A�D�7�HV�fD������AQ;�ڏ�i�5ZK='����� �j�7��� �|�����UԦ�ل���ZY��=���}DUg�}�F�N���G+��t�����=�a�Tk)M�	O�4U����ne��yod0t���0^�|��?����jn���s�Ռ+�W�ԣj%�_ܨ_�b�Ǝ;A#F�JYJ�YU�4S`��r=.��)vְ����4����d���w�}�*w�-o��养ao�=� K�}l+��聾�0Q�'_X���_�����8�Q�G��jQ��ujj��UW\�amݒ	?�Z˾]���
5��-1�;T��OC��Ax��5Z������̪���1W.v��+��ھ���N��ܤ(�re�)�lP�R
;k�����p���S��?N�ʌ�k����o@�}��ڊ�	'2G$E��]Oe�A��(	��q����c���	B����T�յQ���RIjWt���]/<�^s�}Z�0�j�b b@�>�O��q��Z��S!�|H{(�Ϣ����Z�i��.��.�{�ijlH�ɫU2l���SU���^�;���K�P}#�L�Qq��6�U�>X <w���M&�;��S؄w&q@�^�r\_m�?8�b�����*�B�����+�iR:9J��Sc�p�j�&߽�iS��رG���C�O�@=m9�UkW�GV��!ky0�Imm%TV��h�v54���o?M�����&�"��ެ�z</!a����Ef�3G`t�6�[����&��:l_
�6�P��������c����'�DU�D2�B��5�kUw�08�F�*I��Y��H�bHN���X/6=d�ؗox���V�����];b��Ez��G�(ה�+9�J��	Gf\*Ѣ���&s�Z�[U��C"V!_	)�6E���PwQ�cn_DZ�c��L&��3g�����}Q{y���RQ�QwL����C<���ŀ��.��xa�I9lj��m�`�d�lZ_�(4Q��0��,���5hh�	Ke%�)M�6Kcǎ|� \���9b_�١{�{	�/[]�rc��Z���
ʦ��64��O�y�pr�a�XcsV�JU�JZ�dF���1~86�ٲ�������5@��s�̹aPA�^Em��ƞ�I�L2�L��</�&5TC� �ɐ�P��o�+�;x�I!s�d��x@~;��Kg�8l�b����f�~�xPU��������[�D8K��̏�C[7n���w����jZ�jc�u�$`U��-;c�<����b�	�\{���^�������*��C�Ր��!#JE�4�T-ըc�9Aox�[�/���w���Q�=��!i�#�N��3ژ�$V�)��u���%��9B��;l�����z�	�wY��Xs�1���Y�={��&MZ�'�m��	7���Q��>z@�vR�Г`��T�j�j��/�Ԙm
v(�BH��3��������s���:Β3�v�˲c����]?���7[-M�ri_���/&�eIԣ��uИѪ�s!d-�j�ꕝ��;U.7���3�1���)��פq�C�{2��ݟ$�w ���Z��Q%*y�SE���t�{�PKK*�(���`޺5����a'�R1���ȐmZS1wg�1��/~1��Lc�5���ט��Ǽ�{�����=�'��=�s^9������9(F��l^op  ��ٳg�8� <fÆ��ʹI�b.TQ��O�TT��U0ឞ|p�F��|�^.!I�����`r�9��zI��d��C���Y�X��ls���F]uլ���	����Z�ڇ�4rTZ��F�#_]Z����}D[�$U�5�k��ڛ�\��1�����O%�`fL��l�j�_����˦{t���5u��*;B��D�U�JV��m�-*����ԔN�����ZNJ��u�� ���BJR�<x�8��} n���w�뚓K�� �WٜK�`�Sٍ�c �[:ǳ�cP�R��R��x��M�8��=y�d��|����S�7M�6�m8Ԏ�]Y���*�dGӱ��%U��=q���t�P*�S�3f��k    IDAT�6iX�,y���Ջ\���Z���g͚����3`�����n��'���I��q�^wp��wvj�҂.��fuw��Zk
*�	��P:��VJ[ޓ7t��	�q�=�ϪV:�ؘ׽snԥ��T2Q��=�\������c4|䡡VwSӨ����H��|�+�O�	�1��l�%m����:+lr>XCUF���!���� (�&x.�p�����JYj��fJ��ZĤ_���a�fV�v�̘�+�J%�L>����4� <f���M��IM쬑/&�А���V5�4��'��N� �@~��0A�ri��v �E�@�)=���?��E,%8�=,���6wxGf3c�-���؛8b�QJ)ו�,{��t��g��NVk�0-[ܩ�fݦM��� \�ԩ�â�y�:d���+C��	�W�Y���>��6���{�����V�����>���UwwR���7:�ȉ�犪���S2I�r J`U��Ļ�Pj���
PdU�R��}�[21������� �ls��U`|�ƦL�(\�l����2����N�j�
?y����t��n�Y�	{�mG�oZ3���cgQʒ퍊ł�M�)��]��rZ�	S�޻�� W;�EP|:�DA�z�O>�d d�f��jh��m2�T��v���W^yE=@<�x��� kI�[���KK���Ԣ���7:���Ӣ�o��iׅz�;@xGQ�T�h�8�����K:wH���K�X�D�y���m5"������s�Yڶe���S����ZZ�wާ716�0cd��u�H�����  l����/�2�l�.��5��~0�x ��am�q~���N��g� �"�`��^���f�@�� ��`���7���~����^�ʃ>��Ae��m��7�t�H(IC�I��]��&�]�>G�-[��q�lH��C`T8�cMf�(l�6�c��^����4/�v�P��P��[��V�F���"Dvr�:ur�vI�`}fI�ۺ4w��Z��Eez������3V[�t��SU(4�"�	�{�	_��L8קþώo���=q���?J`o
��¼]0�a�6iԨ�n��Z]p��ܾ]w�u���!�����Ə���C��r����|T�/�~������3���g�s�'?�I��:ʁ�������^q-r�6N9��ٟ�Y���e˖ ���`��s��ζiv�`�
̨�<�LX�C�= �H$���'>q�����7to ��ܦbG^�v�ο��=f�^��"�Z����P2�A(�Lh�p1`�!��ݖ���ǵл���`� ��t����p����aՠe{CM6�+��<��CT�@ǖ-���}J���Ot��-z��������/,ѕ�nPG7 gBhM��p/��,�K����N�?E���m��u����Z�r�.�B ᖖ�f���f̸@=]ݺ�������:\7}�M:�4u�t+�a�	".=����6�\����
@���؟P@�`[2�U�\o�����??`&-�9:�@�U�#��3��6p�o~���S/�+'��'|��[���8?�u㉙lJM�-*l���<C���4����Z�z�:;��	@"0���y{Z�����#
+��1� .����f�N�%aI��,0i>f�ZL3g���,�ӯZP��Mw�}�zz6h����ʫ.R���z�՚:�usD�pR�DF��my�8%SDGTT��ل�h���x�D䭵c�ks;gm�w*�\d;6�Hj�kCk+W���gU
ݡ��=��W��|���o���-�'���l��#�Go�t���J�e��2��0vWp��N~��O"Q�!e�(+p
��7�b���WVӧ�v�N>��p� dmN�M�.���:̥�.~�r��`�t0�(���N��<o޼[�&<b������]ԝ�.�l�|���/~���\�� ��h��.�(<���Tl@����~W��կ�0m.0pp/<�쪊M����Z�e�8�aq��;k8��w^�d���o_�!�������MU�	�\֡)�?���&U�TQK�p�@��{��a�)6�;J��1�����"�����|ò��=��(�L�1�Z�?I� �l�r=���Ky��U���/{�e)QYL�w/lҢ7�u��S۰����Cj��ke%��Q'P�	������}V˄��{K��r=�~�<s�k��N�0hB�p�a�4�3�5p��
��/|�g�������o;���
sD*���}��w렂0!jlX�`��'�+EU�5�~̡�����m���_�,DX�,&L��g�5�uv	�H�8r��^�9���P}��![&	���/gZ��bc|l�Ahl���}��f�;c����9"��L����ש��M+�nׅB�E55�L�P;3J*�[O�7����ncfj�J;�vV����WVT|�跗S�����u�ܟ&�P[^��KC5�	ko��=KS���&Xn�r�mڶ������{�3�bK�L��(/W��W׀����0����-�?�;wn����W�vj'� e~c&��=���e�L�6-��f��0�AI���9��7�������L��G[X�s'�Kj�Z9�J}y�A�����ױ��-�Z��;Q3g^��|�b�k�7�~����+* ᥮�6tA�����da�x>R;� ��.�(�{�����6D� 8K^ ,!��$��}�{Ò;���	R�J�Q6-�z��mXV�|I+�n��om��S/e��׉�6u�ƍ=��9� ؄�|�q��+L7���)F�x����7d��p:�$���;���>]��i?���I�$$kZ�j�>:_���F���_���91���
#�+�ʹG�\���L�;bya���as&,��/�g��v�K.�$��(�M��ډ'���ް�x�A� T�;�j�S܇U;�8�29�����=�d�9�;_��v}f���D� |��'��ߣ��ڼu�J�r�	�����j�%9N?��p��A�'M�:Jx�w8����s��9�ӷC3���p�eP��=�RHX>x�/���� ����3�UWG��Ŝ��)<]P*1LK��UCK[HJ񌡨�� �
	��W˄��m6�2���"!N��>�]6Vf�S���
����r�I�^d����	>Ԗ�_�k���{X�BV�ZE�N����o�ӓ+��Cޠ�O����R��U�Pϐ��V�Ř����g�������k � I�*��m�g>��w��L�iچ)@uL���� m̞�1��8D$q˽��1��=��s۠�-�^��ݖ)����E]�����Z�zE0G ¼�����$��!cǍ3T��a�,3(t����2�����-\^�C����͂����aN�EQ/��H���PH$��A�Q�@TG�
�j��ɢ*�h�:Τ��I4�^��L�]~����'���z�:Q%����8+XA`
r.���1+����P�'	�A��%+^�#_���ڕĴPٮD�:UjUe����:b�jic�܆����)��T��ѕӜ��(+��0q�_}��!B��9��SO� �c�k��� p�;S�8c"�i�c��ۨ��<�Wp����q��3��
�ͪ�w��={�-�
�0�Q�V-l�&aFx?J�_>C�-��~���X��P@x�ĉ !a�Ȅ4�S��8?��9����`� ���Z�[Y#P/�]t�!qQq�Hl�@�uf\Q�RԢſז���I���H
xHM�����J� \Ӕ�3��Ã �������~����]B�V>V4f��ӡ�(7!���q��4����ڐ�Axպ���IU�傚�j��u'X�Y�L�&L���*���9�&\VR�>s ����ς��9⪫�
�"A�0����>�g�� <s\�0O=���Kd[3`��ò��y�
@�{::\���b�zI�O�}�݃�#7�\0J���{:��ԪCF����J��.���.؄q��@v��4��q{����YN����l%�&�%�� Ll<�=�%��
�հ���̆�X�����|n�~����ٱ-���
��4;,zi�jlł�!U7GL���^N+E��^�1'-O��񋱩Þ\;�,[�}���^ �d���V�3^S����l�X�f�}d��]R[S�ڇ�Ԑ�&��Ҫ�����>H�}�:�����@��WQ��	��:v��7懛o�9���8��l�Lw����50���
��|�+�r�����(!�S��p9n;4�`�&�����L�"�&�V�~�{�yP�	S�}����O���H�5F��ݺ��[B����%55�v��O%��a�6Nl,��=��H������;��܀V�		AЀ5�<0;��0d�H�6Q~c�L���jG�T
�Aw�>���*�rJe�J%�ܯW�{�B��I�T�M��d�: �y�;�#����8j3[�G3#?�o���f�^p�|lj�o��6d�(0;��"��0#��]���-�J���%����0bs�����Ǳ؁h��a�~|��!�����'c�o�e�p��WHV�nw�3���{�zEc�eD[�N$`~���s8�=��8}�m�A8��Ǟ�O�?/�}̠�7���dM+V���?�\G�=x����<]|񟅚�L�
��R�vmڜS��c�=��R�=�ݳì�L�����7����I�/D"Z��<���{�a���+��2� �I���	�x���L���yLÜ�aA8�o,��p:�~��{��Ƞ�1��Ft�_���v2���������N:F���i�˛T��sw�iϧ�;�&�'8��d b�AS�>Oh���_l�a �����*)q4��>8�x�Ax�ῨJu�F�H�o8D6����Y%z�5e�5�盂3���$l�퍨'����%�`�������	I�\�;u9xI'��~����'��<ϓ؃� ��������!;?׬����:l��\e�fE�wo�j��~��ab��z��������4էhl#7�������0�8��Jn�{B�
.vj���2�ǲ1X��v�ڔ��ξ��&������^���g��n��ݯ�]�A8����ݥ�l�M7O�ԩTQc�5dҊU�U(��N��(-u�&����=F�.�>�\sM`�8�*�[�2�����o�'Vӄ��^����&�6K �=��9��Y�C���>�{s�p*��ڽ��{Ӡ��ȭ�6�t���ܐ��O��:����i�Q�!��~�֯����^BG~tfANU�0�J�޿���&����� �����n#�'��3��L?!z ��z����|�T��%U��o���ƌi�{.<C�-���V,�Ԍ�7��3�J�Y� �鐬1n�X�ӕ`SN�2�k�>sG/H8���qW}�9^5�@h6䕀��`&�I�Ak��{�fñ��@36+<4?�7@���i{2h�1ӴYē�>���ǌ���d�x�?Ã����m��=��$���f� �^_���&O|'�� �qj��L�tr?ڱ���឴��oF��gE�1l`������"�?׫�6� �Y2�e+Vh��_P>ץ���u��v��J%kھ�����J=��M8���%�J7dU,u�S�EdU}{4�.ή�����#��E88
���г����c.��� �ؓ�+�>���w��x����&L;�+˲w�� �9s�|h�A�mÊ����I�R>�Ne'�	�x��B�U+VkѢ�B�bVeA����d<� )��x;��^f�)��{�qR�@h3#�|�|�p���\G��N�Ɋ��-�}�Mںm�.��}�P*����AS'_�Rq��զ�-'�5u��^.�F��pn%l�֎R@�xbz¡L�rI��X�<�e�cv��;E܊�l��f�?�gGGxBs-��خ��������0:�ȸ�eO ���cFƳc`5�5Hr//�<.��v���\�UV�0��0�Y&6�+��9�g3٘�ǀ��C�����y�N(B&1��qR�MQVj;Sd|O]��c��(�X	����7�Y+���.ї��E康����;��5����ݟ�>����6���;u�o�鰠.W�\K)Q��Q��`�a�q�	s����� D�^�+p��j�z�������I#��3���๏A�d�c��ް���|�+�1�|Md��j �{�w�AxĖ�G�J'���)jGx����z���j��	ڴiK��X�[��n�@a��	@�{l+[3{�mz�'OA��9္1Q<�< "�)N=��}���i��c�|�����sp���?������߭�{�3K��U����9������ՠ�U��kRO@�(^@�l�p�h�P�|>������sO��0P<)~����;6�&���`�b��1�`�2-	�=/���6��|h�%��Y%�4�q�������+f�1��;���.blvn6�d�-�U�Q۞m���� ����l�1�s�e+�X�Ǭ�J�כ��m{��?~���to�0�{i�b=����J�iB�c�.��L�x�+}����<\��>W�&�j-�r%/��Jg�D��)��i;~�O}�S�= {�>x@������n<_p�"#c��Am��q�U�My�����}�k}�����d20��	صaarۦ��!j՞��U����9g�+쬁p0�tҚ� ��a9F� F���G��أ� ��3L�a ��uυ��	�e��}ܽS&�H�Еל{n����<8�?q�N9��\�E�ϸ^]]��R�0�z����`U��8ᘭ�^�!����><�]��s��ؽ�I΋Ɔk扣�`�g![��#�0}˃ev��1��ywț��0 t*Ê�u=|-�=<�hǸ'�N��`r�ެrP4g<�Q{�N�dblfMi��oȄ���p<�|�mA���@l;d��o��(װra;|	y1��o@�,�y�6u��ܗ��/m�r���ݦ]�*l��6���KȌ�D_9��pQr���h�s���^5�AZ�)�	/]�D_y��ڼq�:�A��1K_r��nަ믿M�^ت<R��:��	jjlS��W-ݣb1��T�T�;�c�W���r3�3�hcҀ���`EO�\ܝ��=8�Y!#gV|�Ƶ�
�W�}������J�8��MSƠ}�8��6MjimJ��A=�l6�|�G�R^��mz�����x>�T��0����[�D��v
�U0�04��ٌ�k�[x+^��`�;�J����V-Z�s��-#���V�;�`-]�AS�_��δ*U��l�Y�t%d�%zkg�� ��b��&K&�MۘD '��53a\����X�Vf"�6@@��&#�8�}l�o�c�e@��� �k1<���J�����asO�E��,y�|��2�20�7?���L��9^�܋PĘ���'�0�xc��!��u��3q�iE;��ל�In`c�"s+2���Y�Z�f�~�����O����˸�Lm�9!� x  &;r����f���`O�#<�c��2`�{�����{�a��J�+���/�1mݼY�����g���g���C�7��S��TÆ�;�Oo{L�W�T�+�P�,YI�o�p��#���{�+f�?Bvf�V&��.�@lvd��EE5�-�I(`wG��G3o�s3�W��
3����aЙ0�a����*I�9loT��U͔�ΦT.��\*�
��&f��P��섁��!����N,x��`�R�����6U�.>3���F3�@��9o1ס��Y��˺⪋5��B��U��1�P��ZkP��P�rf�m9�
gP�>�cS/����D����xU1���ٖeM��FN0 �6@��D�0�,E �AD�p�m�n��&�FG���w�sv�= 	���� ���$���0(�e��;�0��m����?rR    IDAT� �.5�$@6�H�#�8����D��y�| 2���(@�〓MA�=��g,�8�������_d�,Q���x��w�Mڏ�b����}u�
�!}8��2Gބf��b��ܠD+�FI ��I3n�r��(e���嘕;�2xG�p1���|}��|ɲ���Ǿ������G?6C�/;7���������Rg������c���X�E�=�JT����:���y睁�!8"���0����u�Y�>�!3�nPzȜ1땵��e�x���/��(���J���;w��wܚ=��.�7"Dm�5ZK=')QM��= L	�r�j*��s��t���C�����W���IOL�����}�{�+
�Qs}MlɽA�>���x���0�W����t�k�J�lo���.�x�&L�d��&�t2!�=~�{�K��#a�01� L@��pfr1i�����a�ʀ�=��P���z@���I���	���c�� l6��� Y �s̑h���1 �`E�\�5v(a@�~�=?����o�&�p��$�� 5�gs��0`À KD����r$%� ��XI�=�N����
��K{9ӌ��� "
�����;mQ�\K���w��><��slR���{������	#o���j�%��! >���ڦ������ %B�b��W�����0��	�^�F=�9U��P��;��%�OWc6
�,}iS����o9N��c�N��L֓z�+��z�I �E��<�9�E���>��I�.�߻����~;�/$��܏�?��>�����tz���8�L������}�'+QM�)��� ��Hk3/�c��߱���	 <ӶI����&<Px�[��%)٥C�t������s�\�~��m*�S�8Κt�%S�Ru��;�^F�O�τ��g�2alo�\��Ť�@���yLT&�w ,��e��4|�? �hh� �0T 9�,�̓���n���И��;u}W��r��Afk<&L;�:�-}x +,f<@啓��PZV�6#01Q��s�o�t9x@(7�%���\�yȁ������� ������hh��=q3}����N����ʂsQ��$����F�|�c���W�[���{�3s���y���<�N��������Z�2��� "]�s�ua5�ɒ�ߣ��1��Z�f��ŴZ�G���$��)�TO�g�#Ko��1�)+��aj����x�m������[1 ��}����������9��`mM����- ��=��5�����@U�*=��ڤ�LM-�xZ7��Ѻ�=��޿UWGU�23�P�d��u���J&�}��uڶ�6j�E��<�}g�0������1�cخ�� Y���f�_& ��x���ȅ{���]Lfl���
R��"��59�`E�����1{uH�'6���)}`"��@�z��cF�@?m�� �d�� ��}z�8����N
Ϡ��"`�N� ��?�����x��ov~�^0_�L O�0p���C� 6ރK�"G���PJ���D����w���|'�ŃLQ�(&@�U�G���x������A��B��Y�)�}r�(VS<F�����A��3�/_@�1�R��w�:�4���Q����˵�2�[�U��������>���t�Wʴ�Ǥ�v���-�ܰ"�jثgcW��A>^M�'�ƠD"��x���{��?�=}x�������7�o|yA[���;c��t=: ���K�8|� eM��������G{���L���e��FtC�ح���GZ�jE �r�#T�K&��Ғujn�\��i*ժ�L�,LB�t���m�"G��
/ �2��ق�2Y��a��b�9
 `��Ra;aW�B~LP��L@�8�Cl�+���x �XI�T /�`�8�X"�	@�vp-  �rm��.�o�\ c p�]�`6�➀�}(���>� O��p-��<�L
�8�@�D! s�N����(-��= |��ʓ�Se�/rfL�f�N}��<���Q<�����E?�/Ǒ?�@��q�, �ǽ�@�PĘE����ȇ{�V�y()�j��1���x�L8U��W�s=�J����4���?�!�)�F56��ط���y} a�aja��w�.#[V�����$=�-�=���������|��0�o����W �9b@�p̄-�X(ql�;��`�'��.�53��¬���M�Z����,VO��`#.�XK�VmU2ݢd�Q=łҙ������:z^^R�+�/��b"���y�g��� jdò�A�#��a1�3a�,���d�������^v�"����y�,���4��1�Ñ6�7� ��`Ұl��؃]� F&|O;x>��P"+'� Z��A>�>0=;!�5�{1�A��N��L������	
��<��� ��1�hE�;�g�F��=�����M ��G~8�������v:���
�˸�Ǭ���V,���&���7a���٫f©������W��^SK�Q���U5f����c����C_�lC����+W��)rʦ�;~���66��fKc��{��,����8a[q�����nG����>���'��<ۥc.b�;a�	;��>Y�(�X��,�=i�@�Q��9��5[l�B�U����K�
�'S�+�)6m�-J(�|�T���C� �ђ�/M���T���d��H��l��fb���m�LjX8���o�0N�Cc�����M�q�	� ���
L`'4�&�X�k���8 N� R�t����㏶�0a��&;���P�PnY�6Y�{� p�M�<��w���:~����y> �G�0\��=`�0x�J�N>��c<����L �D��6�˱�$ Y E�B�M��6�/���N�y������$��߀=�����3pl"_��&.�g�=9�ӤdwsowLx��EZ��/�g[U�[ڔ�^�D"��l���V+��c�S&۬D�ݐɈ�nM�R�~
�a��g�8<�]�a ��@H����ڑL&�}���_�'g��5Llnp�t��}a�@�N[� c��Db��B���*�.���׆�W.�`�-R�M�>�LI��
�dB	�K/��	&*��Q�x ��0&'툵:@����6:6�D�c@�L�
83��d� u{G0��� �mj�m��^  �( � m����Y���B��m��eN;`��
����W#V�<`�9,�9F���=����8���;# �6���,w�#'�8������w`�7� � �ڶh34���_�k@���1����]�lA�]L'� xw��w�8oLP����L�h2�{s���=a�ƴ�-�w�wC_ c��M�3C�v혫i��z�G��Y
~��ڪa�KJJ��J%[՝��w�Kc��J-��
�j,��|h?�/+{���x��Zy��Y��g��a_o"��&�zd�Θ�>��^^�Z��it 3aw¬�,ƃ��owfwygߛ}9 ���Rʒ6��h_��Ɔ���-jmI����ư���Et�-��'�T��Q�]M�K/	f�x�v��ba�LL �� ��9*�la4�0,�kP,�c��!�����9:"L��ɲ���.C����� �a��	 A����j�e�Ov�q-��y�U����jh&ǵ�����h�8�u���9�	���̑��> {�Vڂ����v����z�'�B��.�ȹ��YA 3'��S��>��!|���Uy�p�'�w��5��
�}��(+l���A{h�c����Q&N�F1V��`�׮���#��\�*QN*�����/һ�}�ʤ���%57�M[�U��A�0�*0ߔ*�Bؙ�J��V�N$���V��_&>�3G0c�F�h�O�7q���}ʉ�����M8�>�Z+'H[����D^�t"�	aa�6w��Zd��A,6Q�K	w>v8q��߶+٫
��5kV_��_D����R:��a*W�����M�^�Ӫ���K$5u��!YO0[��j$�ι�3 s�D9�1���Q0#'� 8N&�3z8Ppvru(��ISbr��F������@�k�T�}�г�Ӗw��A�w�o�D����>�
��(�X����l�ٽ��x2�o+����J7^aœ<fJÞ��<1��m�W��4��� ��noq���w'�px�ɔ/["�Ւ��N͞}�f�|w����0L�B�::ڴ���̳��z�I�럶ܿm�M�(J��Ϗ�W�摝�~_~W1�M\�E�<_8���=�ұ�7[��7	QTs����W
$k$ʥ��eBD�!c{h��D��~��,�����w�b���$/ `qzk��⥃Y@�]{�}!j��j%�[����[��z����Mo�|��߽�^׾�c��ȆR�,���:uZ��T7��?;���+�y�Xi��/��������7��A.�,��c�B^^��)�tt ���q�Iag�.�R/+�|1 �n����w�;c.���o+���p�T�190��0�K,�e߳���e�6�N�1���_�|��+�݁���k���/H�����{�L͸�\%Sm�Э��vc�KG�=Q�v���X.)��(A��2���!��7��x|���v�ج�I��q��oכ���c"bR�Xi�!?�Ǧ3f�i�`\I�Rߜ7o�5Nػ-7�;��\����p�݉������f� �M1S�Ϗ'M�<��3 ���ۖc���`iG=a�t&�c����G>r�
�����t��h��az��՚5����ި��)M�2]G�K(����5Vvd�ē�6�Y�Ď�ͼ�8�.vDY~��Ks�-2`I����Vlv*�go�Ҳ-��F�d�f�?{g@П���Z���u���?>޷�U�p�~�ցd�������$ f�Ⱥ�.fx�] x�X�N�>��s��Қ�w����g+�N�����>�����ܷ��}�4�t�
ee���)��L��vY;��äͲ�j���z0�8z��m�G^�7����Y�Wp�o�m'�Y3�2�4t�p�o9p��έ��)���90�r��R��J��'qƘm;4par�`��U�i8`�q')xpƬ!��v,��h:�~�q�мf̘�g�'E ��T*���>���~���М�7���&jŲM�r�z�[T���� l��[+m�i��;�ENQ�ض�	�d���,������5��<�cVX0 �M�K���1V�����+v������x�����{P���3���{�t���9�+6������;�>0��uv��l�*=�p��][�>��;f_�K.9C������}���i��7�;�ao�r��a�M*�����r)v\�v�j�oV���@إO�`��ybY1�#�1��<��.��0��8̔k�)1�ơ7op3���ǎ�qՂ�bω�0�R�+J4�B����`� \Xv�� `zY@�܎�t�[&���2O"��]����G���Y.��eĪ��y����Թ�C��{���(� ������g��eK7�]��T�֮j��n��}L�� �΀�ϵ�����x��) ��o�a����l�f��2�HM��g'�#C�K=��\|����"�������s�q�������̹�;���|cv�/e�kNh�������ڦ��U�5{�.��Lm޴I7}�.=��f�s�n��^�w�2#���Xަ�Ɣ�lWQ�9�CD��x��ؔ��31�`�6�`���'59���qm�o\ɐ��T���
ګ�}
��^wۑ�����jI�".������	�1w��G�XK@�Ѩ�P���Ll�r�=���6Qx��tU��Fx�/����ĽB���#x��Ȅ�ӧ�4:��:+��f�}���K1�@}�ԡ��ŋ�k��7����0*(�p�c.TQ�];�\n����M{y����P.��?Nրh`�
��7����6���r]7!vJ�m[C�.�3���.fb��eg�����
��;s,�a�1��@�1���،gv��0�=y�@�����X�Ǿ�@=�4|XBw�}��N=G۶l�'?��?O�B���ןt�&w�����.���T�ϟ�9��V�g�uV�%|��I:�EH�&���*~�6]��
���́6IX������+�x�o
��p��/��?�V:�P̉>�m!:"W�Vsk��1N�&�4������fR#DK.'.�j� ��kw`���s���XQH�#�"�ŕ��������xІ	V+�\���wݬ\n�.�r����^���j��k�+`nQ�<u��7^rPB������`��c>�D�����˯���8^�}�c}_~�
������]:ۋmZ��$��企�lo�lw���-�8raW�tO��33���	{��}q�.A8Y��K5�#*�t�m�t��4m��x<�̏�K���ϫXn�M�Cc�zk��L$ECM�|��ɺc��6�c����o㋽�\�H!| 4c�ӟ�t�W����^�r.�?ĥ�L?��+Lp
�φ(��'��g3o9�5M"&���y���e/�W
'����\S��.��l�1�Mԉo����B3)�1 �d�1��7��v!t��Ht�����������,x��~z��E(������}:ċ���{lی ��u�?����z���*��V�\֦E]p����;kXKk��+u�Q�ao!}�^Lxg`3[�#l�I��[���(�3��Td{q��7��F9:���!�A�n��b�pVK����_A8fJ���f�x��&�3>�M��?�Y�'����p�utDM�V.����/��-�[o�����U[K�:�KZ�l����s:f�)�d����^B�j!�Q�^g#�	�NoBxΛ7/�ѯ��}�帆﮾��0���6[G�x�ސ-I=בI�8Nn�w?����0�܀2��duȜ���w�sO�{ｃ[�}��|��Mk���r`#J���:n�&O�4�5��z�kO\:n��@3]w�F���R�� D��sx	`
�E{}�������*0�_��^�Č���5aK�n�uޑl�7(ky5d����!�Ӷ�5�6�Ce��/m��_�B�AU�Bմ��M�RG�=��~��� ���۫ /�̈��_�r1+f���Px1�s�u.C�����D�_��#ݛ��}![O|�W�Ǡ:��&3Ƹύ��Y2߹nn�t�K��I�q����jǽ����@���Ym��HT�l�-\���;�jx[Vw�y�&O~��U|ERcS�:��Z���9٘!�t&2n�[��l9JYƊͅ�0E�w�y�}B*,w�����׾D�P����c�g�F���1�l�u}�wl� �7���T~��D��H$�Ycp���Gm^;����6��ՊԚn�ȑ#t����[�<\���9mܸ9h :e��
B�|BM��}���q�&�Ɖ��6��\�i�L.l������~��9T���k=>����=��Y+(��Ѷ��LKɜ2e5-_�]���W�6��%K�ӧ\�qc�V:�Pg�$lP�g'!j�����p��
�ūgG1m{���I��]��w���cQ����������TzE�?�0fz1 ǡ��x��α�|g��ګ%?�J!Ί����
�^��db�;�=sĪ%z싏*�ա�mM�|��:��w(�%�?���(�fK�����$�4U�i��0G�2��~�0'xS Lv0YL 8�#�3\��?��`^��	�ZVvA�ۤy�vx��5ϣĀ�R��3�J}u�w[�GoY7�9���D�sò���t����굫�Ң%!D�F0�A9f�Ih1j`�y�駃��n�Pb���g�}v�� S�?�q_	ź)�\��2�X    IDAT@9m&Y`;4z�ZT�ܭ~�_�e��P��L�j%�Jy�֯�R2դr��Z���UM�2K���t2[<�w�;[�ƀ�h�]��}����U�d�oX���۹����-�����@pꩦ�o�ݫ�	�fY��������
�����n���1��Nc6(�~|3�o�
����_Z�HO>�
�|�H8��U�ښU�w���g�E��S4z��T����O��a�k�U��W��v>[a�'<�|�M�b �܀�9+�&H��"Q��b�\l�3�����e��C&|Q����:��>��~ �<\�����}���!j�L�=�#�V�P����r��k+`�%ځAb�o6��/ɻ1���л��J`u�%xY�J�_=N0�jQ�D i@��E�=�b�SJ��[TcC��96m	EH�	v��	�w����
���O���`��'
�=�<���v�>|G�aL^A��v�mF�Ն�ӫ�����A�w��]k��� ��x0���!�mG�kT�p�!ż��n��l���۱+Ξ�#��Z������խ�tF5̉Y�6�R�*j�*V:^�)�*I�%=�L@���U�Ʌ�K��o��P��F�]�>�7laFr��3�-k0�)l��X��vk��W1��躐�ìA(�O>
C�,V�U@��s�νip7�����#7���R�>&�9��чh֬+�S����j����`�A�F4ڱu| �l�6��BC�N��`8��s�	ڎplϘ%0e0�|� �y���A�~~�ew��\T������B��v%��'WS&�Q!׬tf��h��.�eM�
c��1s��s�*��Tcd�l{��cgVe��5��U1��펾��ڸ7���L�;���<ۀ3_��ݫ}��n,�X�Y9%66),��8����O ���Ήw�v��/b������x���{��0s+V걅_R��G�DM��6e3 k��ʨ��j�����<\�dJ�f���3&j�@n.gi�1��v�m_(|�s,��{�E�k E�E&&0�|�6��{G>�]��^��^�3��Z����o}K�j}�@8�zjޜ�T&Nx��� al�8�ƿy����*=����_P��ҫ��p�1`�DZ�P�`ԟ5X8;/��'��h;�'�k��&����%�k�n��>�9�X��oK�͋E�|x�9�C0�Z5�bn�~��h˖5��ra��d�I�|��.ݢ$�Oq�%s�97}�e7�(��^		u����&>>��g�"J;]��Yml汼͢ݦxij��g]�j�h�nWv���y��f�՞cZ��#O Z��Vef��x�j���6  Kq���{��7�
Kwf�**fz�{�$o-_�Z_����uu*�(���M5�;aӃb1����\�g5�ua���sy0}_Q�|�P�����sa�l.K�m��"?�l�!�L���k�{0�T�՜�1�����J��^�rh��v�S�$��ٱZͤ�_���9��[�='��|�	�8�m�2e�~�_?Һ���UQ��8�H��e;q"6	`�A���Ʉ��B������ H�~�,� �ܹs������߅R�/����c�?���h��$s:`L��s�C!�l��_آ�n{@[6W��XJUKV4m��z��`JKb	�e��}���~�~�V`\g���o�|�X=�|����	���N�ݱս��1�}�l+�x%�@�(��\��8��e��M6Sp�:�*���}ضH�0s[��"���2�\}϶a�Ǹ�� c�s�&�zD�����]�)�]�A=���/{g�wU���]g�Lv�UYٷV�E4 	���
QDY�E����Z�B
T�.�V�\�hA\ؗ���$$�}���~�?�p�w&�dk�:וk2��_�y�s��~���tw���m�矡Y'q�`?�g��Ʃ����^R=[��|~�����L2��eW9��,ކ�x#&]�5!��"���� ��c����
pSmyĆ�棵LL���B���;{��%#S�j��$��h4���}W\�ы�����;c�m�۬Yvg{��P�lX���	'�E<|�֭_�j�2��V�a�µ_�:K�P@��\�a���p Z,�����ٳ����a�qx�OX8B(�]���ج��~��5( RR����T�s��պ�y�K��~����������k�<�0 <C�75����k̪���1b3d����1���f�1���m�ɏ���A؆(��l�l�F�G�4p,��F&8%Ly��d� Ą�p�Q�b`Hb�f��6��*� |��q�et���@��������>�a�8��%r�a{fɳ���w�&�e����B��z���n囊�h�:�2Z��/�`�U���Ԩ'��S��L�a�q_�Q�>餓��#E��z�	c+�Py;��
�L��0(�
��, ���W�}�,a�p��kO`��+W=��Q#&|͂�;찱;ވ>۬}a��Ca���3�x�	����*0a�#PBvj�v�Q"��'��}��G��k_��`�m������ �2�����;/�7HUÅ3���s/ ���q�W(���{nծ����9G�e\����^X%�z�T)OR����蜹��mӶ�1��%~5]�6�R3��و��04oAgl1�\��צB�N(�3��C�(��PF���CHG2�i���|�.�B� @�>3�a�� `�=6�iO�@��a#������
8����=ٸ�~���"��T^0�]s-[Ӳ��ۿ�j�&�gt��wi�i'h\���ݫ�>�L?��ot�NҤ�;)6����2�����Q~ I��:�������pe
HiE�+Ű���½������� n�̡d�_�	��˹�������g�;��5�S��V�\��]{��c^�rʺ�'�ˇQ;�z��춗�<�=��
����z�,�a�q-����\�b(
�b/`�-���=��&fl��k�b�$V�1(9+�>�Ɩ9v�`u�����2����e�]�re��~���я�7��=ۥYo;G��dU9�)+�9s� ᰅ.)쾙y�[���� oW�3kq��<q7�.�38b*.�v�7��"
rT<�_���/ڋ~9�;�}f���"�O� ?���7���'��nﲱ��6h�͌��f��\����������s��v@V\����3?��Q}��E�'�/�×�Ws�Y�J�~���u�u�V&;U�/�V�L�_Ŧ�����BzA�L�~D[b���7�����v�ϥ���'�0ǹ����d��0@�X�zꩃ�`�Ƚ�,��(e26�F2*�q�\�*����Ύ�Ps���c
�u��v��q��ÓڟE��v�駩yBQ���*��I#Q���q1�:��RlmF �hX�?��?�O~�q��!�j!t�q��^��,qA��dל'��]c�� �(uU�L^=�}��k��C?��{�����N;３��J��K��UTU�h� �ʑA�<���A�ƌ2�N���%�ڟX��1�C(7�I�7�.^C`�1a�1ۦM}?�^�H��}mⰾ��Ô�P�d��z�Ā�
�����L@L���sx©\�� .�|�O8�g�p|?���>�)�Pr�ʗ�铱yy
��%O�w���f�����|�9�M�бZ��S��7�S;l��.����^*3�5j*���U�JJ_���46��;��oX�SА�7}���?���&������:+�^3ރu���$���+�c<���8$��n��,�J&i��\������c�S֬^�V�=&�f�u��o����/�Z�R))������U`O,'Dc�}4;��VpPRL��ߞ��f)o~�C�0�0
������0�T؋�,:8���Á0���;�OިG��c�Ol�[.�|bX��~�zzra�rEQ.�}�W.07�Gl��ְ�?�{��� ��xO>@ȏ�c�Jf��b ���+ء�g]yW!F�%9}�=%��c��+K���Ϝ�����9�.p�qh&[�z�ސ�5�VZ�jc�}�Ke� 4���Oq1����\!���I�FhP���I�� ��h�%������jG\~�_�z�ŗ\��=��&N�S�_y�v�c/��P}��W�a`ja{3?1[��#�<*(y��ؿ�����%�I���<�`�@'g͚�@>L5�#��F�^��1�`A.���ųY�C��|�� �7�����pјo�s�k�.����������O�v�q��o�;�����Y/��X���
:�%Y�d+ ���"On�<���qز�\C���?�?Z�h� ��� R ���9w�DҮd�)��:_O?���͘��}��`=�||���=O��#� �`�3��HU�6w��O���X���8����钂C,`��Y�</�{�_�Ťe����=�ዑ�a�3#�k���LPқ�2��.3.o}u{��i<D��Bs���t�<�m֍�:���c�f�2 /����\��szn�
ݵx�*}���.]v�;����^����O�G�L��T]����w��P%��l4 /���,r�&�0?�H�͐7օ c�kƌ
��#���w�uW p��6b0W��3�fԮg3`�o"���cH �9������Y�p�c�S:�_���uDH�md�� 4���o9JG��Z�t�{� �X)�rc%�o[d�8�@���.=�oߏ�8��E9��(��Ua�U�e|�M7�ϓ�yIa��03a�>�eg�������J=����y����?+���V�\��k�aa�Nv1��9M�����#�ir�O�Y�Ȍ	c#135h�l֬8��oJq8�L��w���7��>���9�q7w�~t� l&N�!��Y�S�b`��@a����j�fo����6��9�#m�� �������)�I�ce��ιD/�[:C1᜖/[�;�r���^��Vt��gjC!��������SWW���˴�A�+�e��9� ��I55)���E��ǃ�K�/�����
� w�_���<x`�?���y�I���FF�����t��4�����>#���;���f�s�7^0s�̱ˎ &�Æ�wf6�=��OkK��e:٫v�NG�F��k���\��6���n����R�!�3tP�+�TK;��#�p���*��=��u�-����}H�'O8Y L&N�m�?��{�u�&��Q��)T�7i�ҪN�s��;�Tm��N[&;b��M�[�|%����o:Oxs'���u#�Y��8�O#���I�m�q�5f�CńcY86�g�0��O��z9�K��m����7֛8�����/�F�����\됆C^���q���G�����M`םv1 0p���} ��h�.��p�ւ��+V�+�~I�r���}��Ӗ�<VM�eut�����Z��_S��	S�U���,�ǩQφR�6.��4U��m��c�]j|�f��/�8x�dE�u {�Ћ�>{�t4v����"xl~�z�9k�!���b�.19��d�{��7�o�AxʚUw��&�-���}5��4k}�:��N:�-o���3��E�⣋�披EpD�)=Gp�!:��3�;wnȂ`Cq��|�ɧ�ӟ�tp�H�p+�I�r��0�es� ҡwh�6���ӻ\'e��W�ӏw��9�T&�٬Z&	\͙�A�{)�gQ�:���ູ�	�q{af�N���� h ��w�@g]2�3�t@����e6i����~�C#�g86S�-��Ôx�/~����Mq�3o��
d��q,�m�;��o0C~�g��]j>�����=\u���𙋔6%,�nݚQ�0�E�s�����+�>G�N;^��z����Fmmؘ��5%e���/��T��X�J99�֍�a�.eI���O|�t	9��w�������B����c����c�l��Ϙ�a���Y!�l쩠���F����r����d�)f���RO��CY6�N����k�����;�J��7T �Ӗ����i�v־�N�0��(尢�` �Ap�k����i#f�qY�$��u�[Hb�(6��=�"V���cΓ[�0O�֮c�KY�|M���6�j��N}��VwWC���ҬZ��Sg�����G<����H`�%��t��"�}��w!%��x;퉶��f��JG�'�}L,�cc���ص
,�F`K�{O�7^ȏ�]�!@ ���3���6
���33�o�_g
��.�E�c��$F{ i�0�z�F�s�{�k���X����>o
��b[��1̗ԁ�A�ٌ��|^���e�F(�_�k��x���d�IH!,�LP��I���V4i�����!��d���,+bۤ��xi3&�Z04ȋ�g���%F�c��� �C=4Md�z!�qhgz!_�1��p�����0�_,X�1a�&�_�#̄a� av�UJUm�������w���	a�Pv��k7�OO���"[�j�&�$��L���7�'��d��n��"A�ܩ_�Ǐ���uji&e�'1�f=����8�jU���ե9'�����;}�e�-�?���:-9"_� �d��;2f�G�v㝞�1���=:D�p�ͨ�<Zy�G&6��
&,��o�Hy,#/�!?��b��1Nڊ�a��nב���gB�v�����6�@�#��i�`����y�Á�#O=�yµZ��Ld} '�Kjd8ȳI��6���4~�P��y����F]��a2$�!�D(�Fǲ t٬;G�;r�%B�����i�����'�`E~ ��s������l.�8��
�x��ⅹL&�ʂ��p���f�	s�'�lM`�J�w��p�*I�C���� jf΄$��F�q��V��8�Y�cA{Ų�U�B%�Z�[��U.7)�oQ��S��B�Rk�z�f̜�l8i#Y���{F;����GNL�H��zB���8��8�h�06ncNXw�'���X�F�n�J�C��M`�Lf�D�5XY�&=�3ș�%�IL�Ek@� I��A�n{�6�a�� Mϓ��� �/`��C�m�	���%?�qzz��}�=�\ߡI��U+�(ñaY�T!\פ\�5��q:;�7̽z���0���f�p=��|@�= (�A&��K"��9|�3����f!#dF!3���⸱�o&< ��]s�5�9��~�m��#�c��<�1��Yi�K�"����PP*�:l�	%wƅ]���}V����|��SO����5���W_O.�P�\��+e劍~�s�Nꡪ�T8�O���0<n(#��$wZ��*��s=Gۯx>�	0������*�0ڶ�~����	�X����X��۸=��i�=�x���quH���L(�{7 Y8��3&�K0�a�a���c�����f@x�[Lyi~fٳ�����b�Z��U��J���y�T�*[��n;k���z�31�$�!��/��!/���CQ&�$���ymo	9y+�=a�4��������2r�VlD���=�=�rc��o��׭Y�^�=b8&#LO>[y�+�1���H�z>� ̖�.���0���v���K�A>V�F��J�[?�����g4���<M�d��_�bq��J5�
 <�Wف�ԯv���)!gLw�,�r�b��X����)�Ϫ?���c`L��~k�wS@�w,ް��q���F/�ŋ>gB��8��	n�Π����]_<�u�>�B&�P�<�������;�._�ܨ%�̼v�)6Ȏb�˟5�{zU����o���&�+����/���=�~���q� ��,�}��I=��2����EM�1����X.C��-�{�<��X/N�����j��L���P�1�k�\.��k���1e��׼����7��0[Io�$4 ���%3;���@���Yn<��3:O,Ѐ�������ꓢ�#�F���zC%��S�}D-���>E�>ݡ/����    IDATJ��y�W����5�a�����CHt�3����"p�PL��6�CyE[
�ai�	ב�t�K�c�����0D��`��&k�svv�x	��p��U�gx��Yxy>���x�;�`�}�'��X���W�?��7� ��8cǼ ������M��,��dɬs(���ҥ���۔���ڒ��Kޥc��3�l��H��/��Tn����q��T3�e[�� �/�^aQ�� ��`�l��cꐏA��3 �X;]��}޸C�A�`���M8r�ܿ]s�5�" �V�=�U��1�d�cR�Ó�V4IKv���`�.XZ�ce@x�u�Q@��;Pp��k; �"Ύx��������zVi��NRKKU}�u�x�����is/ToO�JՂ
MI���S�j���+��&�{^�1a�U��� @�:f]6�1��R����s�����>�$�[9V`<��3@ ��������	O ��kv�N��]XK������1R�.���j�T���g"//�J 0l��Y�">̵,���!���{��_B�rZ��y}�/*��Qss����<�:�8�8�F�e'��?��ϭS_9���I��,+�mW���z%�}�=x�v���]�*\����c��A<�D^�C�\���z/�ǀ�^�0y���^�ך<nc���l���]t�n۽����K ��J��Ϻ
���՗\[O�TS�x0cv�'pz���y��E̼�!\����f��ٹ'hF�u��O�-�f��:􈽴��U���:����vMF�ZS�X�f�</l��e9$���M��1 �S��
��-��0>��/v���r�7�o1�<����I����c�����h����z���AO`������ ���y&>�矋T1o � �k?��={y���e ��s aV���qX�g��1>���%�>�&�՞�e�� �r�*�~ۗT��W{[Y��;4��7�ؔQ��^������|Z�F��^��]�ϵ�\��X����~6����#[ד�m��蓳Bb05��`�޲u���!�� Ӎc��t��+
�ۮZyW{�/0a�3I�0��3�cf��'��	Sw�k<��'���v���oTQ3x�%�8C}]r�{��������U�/=' �SOn�;Ϟ���R.	�d�Y�}���"Ȏ0�e<6d�ԯK+��(��`4���c,��cθ�~@hF2�c7�^�3�T[2q��1��粓
0!�ҋ��V��d�� J��H����� ����Ʊy�c����r��llr�E���DV�1X��X�c�5^$%"a��8&�iC�ӳO-ӽwߩr�[���v�	�J�O���[�U������aG�H�}��vI!�I_8���k,��	Wz�ƞw�k���C#q8��3����r1�dan0�0L�l�\O�v����t�A��wbS f&�8��<ǩ&���	��H.���C�/�ȫћ��_��~��������w߽�rEI'�:G}�mR�5T|���'���f��ˊ��qrR�; ;����d'�V�t��bH�hDf�V��P 3b�,�|�&쉵5r�{	y���[�E�����D.�8}�3>�6���͡��A/$�� /y� �]rX4��&%�6�� p�(`� !lݛ�_5�L{�U2�rZ�r����ڰq�&���kߧSN>>��-�����2�膅�=����4��3�'dP4B�D� �Y�Fr,�'��=`���A�u ��M��rp�����.}磌�:oLO�skW��^�ga.�?c&�UR;!m=���غѱ8�.fR�	��|}�J������
<��0�E�;�Zx�U��#�W넒�|�Bx��z��:������)�[��S�N'�r�^7� ֆ2��D�)��L�?�{~6l�9�W�c���C�n�l ��Ӌ�2 |f#�1�.���a��O��X����������C����0;�`�;��da��o&?!<@�����=���;@����p�����l$!E�8mlH}dǨrz���oܫ��U�<��˯�K�4�Xm���/�F��2���?�j��?a�J�^U�%������4��Ĺ�c�A�n�����>�(�XZw�=��c]6��׫����1a�-OzaL�s/G�Y���Asw ��y�o
��~9��-��CV�pލ��x#?�e`]/�s]�n��Z=��O�������ߠ=��K��a��>����ʩ��4��P;��SN���,Ւ����WyQw��^�0X��D+}<�caP�X]���+q4C�#f��9O,_?�e���;E&L���a��S����v<�� U��,�x�Ӽ!�qd�7��4%�IZ&�)��8�J�:�@jZ�g+&!6O�>�\�l����E��|^�ƕt��h֬7���G7��	O���>���w����\PWOg�?C�B!�$���nCb�6q�o8=2�ݔ��a3/��ld��%��t��\�y�r��.\���1-e9����x��r�aÁ0�����]��c�A72�'��C����5�\�x��B���3�v�i/�	�n!1�Z���?z�j�U:�o�g��V�g�u�POOa �{>����C����B��"3�E!t<����d�Z������G��ً�+�|�p����Y�B�	�`FmX,����E���/�]�>��t�� ��<p��ɒ��]�B�qo�u���v�����'ǁ�qg5��|aT��w���s�m��oPss����b�|��d������?ޭ��Ї/�V�f�l�(4)�M�- L�i�6<V��i�I@�8{����vl�z�U̃o/\��}cz�F8����{u:V�'LL�ě5L�T3b3��:0T�'�n�y��<���B�e�|O��pD:&��S��>��oi��:�35uj��{���ɲ�<=b�N"��#V�'�3�z&��11f��&�P�nk@m$�{Dą�o'��<��f��'N.[���]b�.a��a����~r�d�m3�r��a@��7�:�d���=�F�v��]�)� 2� �yƄ#	��|��9D��C
��.yN��M�z��Œ���/u�)Ǉm���=��J=��J��4�����96rp"M���|���a�� �##�����66����8��a;�wa*/�zm���#�s�ܷ������9�~�u���!#�0����
��������B���=1���-O��@`B���cP6X�r�7����8;�q�
ɰR�Q�nפ�vjҋ�*��W[�6z���:�����ʐm��:��5t��yz��
��$=-)$���y,�x��A�1 !�ȴ���X��.��G����?ވ3�V۸C�gs�֦&?�u.�=�V�3�+�b�Q�7Ġ�^F�x����D_��ec
�dl���8LF�_�%|P.�n�;�q�pQ߂����K��2��@�*��زH�khժ����I�r�&L(꣗��S�E�:E�
ji��Ξ��[�J�FA�-����W1?Q�|�*��"���\wi|���3��u�{\�1��I���PQ���qaH�C$�W= �ߢ��A�����M��|��g��eԎ8� ��q5�#��~Ǡp�Ր^cpuz���t����W�bBL�=�0�p�����3�(ꌠ��Y�����7[4O9�A���a�TQ&ӭ^xF�dU�_�b�-Z�lI7��yuvV���T�t�����9� e-I�ګ���|c6ʢ'qa&w� ��cm� 	�2i0Ƹ�^�J�Gb�ǵ%�&�W���'�}<�@X�� �	@;Ǖ~`��k���o�8�.�@�g��u���ʞ!l���dC�>�o��!D|V��Yo�c#~�K!�Ax��%�p������>�zӛ�T�ҝę�ֲͪjm��b�8���a3T���ib�I�=�$�h��6'�5�c0�G6)��qp(Ƭ�G�a����wv�;��s�yޥ�N~q�ɍ��=�]a�!�J�,RԪ��fL����>v�hs\T3$ǁ�������Xx
�s=�q�|��'�|������S��T�{����˘�(G����xw��(mz2�uU+�����]}}T���">�RC�R�::9i�|�lO؜2w��|�5a��$�$[�_�?��qYD����4��e�͌f4rQ���opӃKY�
e#`#k�7�`$wכ,�61��G�"�!�`١�a!l��6sX;��l�� SH��������~y����Z:r���;�YI^�p���"}�Q6TQ[�b�����HU�!7�6�O�m_ԥF&�RoQ�ﰫf��&L����B�����dיK�z��c0b����7��x�	�S�X�d��xa�s�%�����H�Er��k��g�End��0�T@�Z`��{3coj����L&�\8�Lxƅ�m�v����(`^�6�s�zM�BU3^��������>!� �ԧ)�H�Bh6�Bz�:��@3�u��t>��yw�q��������PV~��o�&�0�c�9F���g^v�	�cZi�|��!$�У�>�Ro�����^M?I=]R�i�*UJ5�l_X��{�ٚ6m����X쓣�^�?6`���DQ`�;p���w��h�³�*�(�C"f��-�4@��|4��^ރ�xLlBo,|yK7zM��v`��d�9�� ��3���f `��9 �x<��x����`D�`ڃ�nX<�ט�,}��{:2�#�>�;ݭJ_�*�t��U����q�p|Q.7A�}d*�IS&�yCK�=�s�0�I�tE4�O��	�����a̚����� s��� �k��
+�'�`�]�ݞ��u��`$�4���K8 f,h+����˵�^{ј���,j/��p��b�®{����6�Ӳe+B���h�M�K�@�J"4�]g��5 ľ��m�Q�N8!��}�����gs��fፓ5p�-#�;��#f��3U�to���K����~�Ҫի7j¤mU�g9S$Z@x��P|>O�N�}u�178%(�A���j}�������|� �DcB�v4�Ǡ�c��Z��L�/nͻ�r��8%履�#�it]d���iz�d���M�H��C�`��9o� 0I�7��p����w�6��� �P>r�^.�X'�����%����kɲ't��U�mRS��\�W�ҋ��-�*�m����@esM��	ƫ^�"bF�}�P:Y�\�+��8:��@��tµ��r�[�s�}�7�ac���H,3��ZF�6�`��]�1K�����1�e�Y@��c��_�hۜ"��<N�jV��m:a�����{��?@ؕ��xfE^0�$!4�±���㸕'2�b���s���(�u�]����x�_+������ٸofo1��چ�*�6�_�s�:7vJ�����sEe�mz��U��[U�$i4� <}/��Ձ*jM��R&l�4�dl��3�2X�<�1ak@o�{̬�Έ�7���x�I@0���ۣn�;�>�X0�	�9�H��l	t�z�|a����:˖���?�i Y� �ș�p-2�~�=�;w�0�F�VM�
��f��UH/��?����5�vJ�JI;�8A-�R&�d0��8q;�|���m�}T�'������{�9R[ɰ���y1�~;���81���w������'�3�� ֐5� ����*{��g�l�����³����p�C��[�^��r�o.X��c�SV�^4%S �i��9c�~�5�Z�f��z�i��&�B�*!�3�!�V\��N��� �^���{Ă�"�&9K�$.��<�����o���ͼl�`�����o�)_�R6ӣ	��U-w�����{d�.��@�	��4��>��|~@yY�|��YO�f �ǘ$� ?('���΍�lDc��g��@G�0,���Ys��Ѿ{S���KX��3�&��	�sl֠�.X3���C��i���y �s\�g��\W��0b��;�U��)�#1��K��60�'�zT_���j��j*J�;O�f�\�B�v���ꮄ�����h��ev�����)��2����A��L��+d�gȒ�:�$ ���y>��@,���:gW�5��N��^̴�y>�s �{�'`��Q�V�����r�!��D�6��pso�A�����+�SN����_��~ul������r��s�(��M����(X���ٚ̝o�2���!��8���dG���e�	i_Ҷn)�N�nۢ���ɒ;ث���z��:y�{��פ��j �,���|.�W���dDff+�9ed�����-��a�5�y���5�d,y?���y�=*��h�vS�g�qYЁ�B�K��d3��j��/בֆ�9����@�(I��x�f�qxs0�����s�s�E>/p&��49�Zn��g2";��/Q�>M�ׂ�.Ҽ�OT��Rؚ[����auu���P�S����d�l O�s�v�X!/�
#�#p��=a�#�u�r�l����N
�x3�מxD��.��&����7^�䏐���Z�V���},�xLA��)/>������B1�r��ݷ�U�z�;�b�Z=���b�1~i1��Sh��`k'?v]qP*,44�ů��\���Ș �����Ზ��<I�܊��X� n�У�~����L�)sߢq���j�ji���U�o��j ab�a��K��pD±��@�UL>����B��N���l<]d�c�:���3y�R��}���� ���@!䙢��a������:�݇��aa��88�y.a<FdͶh{0~;B��q ����Hy�=���l���m>�b����/�V����u}貳5{����e���o~L<�f�8R�l���
;�Z!�̚
�E�O��zǜ�l,[���!�����!��v�w�y��w�yg��E1�1�d�<`������_��R�����{'��"]]�֢j�|���^���1�k�/������NJ=h�:�y���%O�t�#�0�!�Kh�]4&�Y�Wym� �\-r��c�y����F� /l��o��E��{b�P�L8��V�z�_=�kt�՗��g�N>�X]����5�G���y���E5��x0�/��9]Ӧ�|XGxɅ{��0�J�Γ�c��;��Ŵ�ٶdru�W��Qy�x�:���nh/`mjG�h�e�r�����β��i`�,�՘�S�(�ü��0�a8.i�-�0a�8���c���N:d�35�����d���Z|םa����U}�w�3���?y@��?j���.�kM�v��բ��%�^V6Ǯ��td������aLa���1�<�G�Kb�,ԓ����O�!ț�8)�5�9��)������Ż��l/�﹖�ID t��3ٺ_��j�|��kn������o���ֈ�5&�Z�hJ�q ��t�̃C8��?�ZK�?'��BH�0�
���;n��P����.��� ��[ɉ��x�A�l�@ ���g�pPZ��������p/��@���(p`x����_.�u�]���zXS��붯��^��nz��:�B�F�\K�u��9�����d�k>ʓ5�I`��} ���zP���Xm̈�DF{-�i��88�?�b<��{<�}�A�߱[�^�L�O�����[��v/��3& O�u�sp~�Cc|�gH�&�5`���x����yq=�0��L�|���-c/�� ��X�hb����V��oUϋ�0���^�N�|ʛ��]�5�������4i����G�����U.OvUF�ZU�BN�P'Y셩k�I����J������Z�#;X��?��p�����xA��~ثpx�ޅ�:��K���݌	�;2��}q���E��W]=L����~h�I�W�9��H�VUԎ8�0�t�,���/�n�ZUJ֓�5X,2|2�����ut
A9�������v�m�s^q�3 �-oyK h,��,>���0g���_�u��9vcE�qa�sl���S��c}�n��:=��o5~RC7�C:��Ѿ�q5    IDAT�uݚ5���4����Z�"'���	�MQshd(F2�Lw����l(��y�E]|��~;��+06��\��㉀m�B��G�V�5}��I�3�aY��x?� 8��6Z�M�v�g���.f�<P%��� ���qȇ��0ۀ�� �2�ŋ�[�+᧟Z��~�N�z7h�Ć.��,�tқ�am�.��=���~�}��_��4S��b}	0��/���<�f]���g��n�A.0�P��s�f, Ɛ1Ǔ�]���3�y��X��;�;9���	��������6!W�AX�b��֔����]~��z��m[�#֯�����P�Y�����ЬYoӯ��־�F}=����D��d�B�,OPB,�58l����ɂa��
�����{  ��Ib��(��t=a�3a/,�)�ro�nXx�~�˟��Cv�?|�Z�v�]�?,�9�H��Y5���
�e�� z@���F�1�RR�g��P�?i��f��<�q���s�ꭝd�N߁�X >c��ǘ�۬�qf���f&���K_gC��5{"�`e=�6
�k�x>���c��aWN��"`0��.�,�9�3�7�^�Mf��K�¥��\sD���"+��a�n��~���+��[յ�M����׼S�g�Ύ�n�����>���t�?�LW��)�Y�(�YQ!�{��Oh�e�¬R����w�;�l�r�3�����_���s`��#L�x6^��+��m����Q�QJ��"�E8��R�T-�͎=����ի�l+��R�QML�p��5K��G~7��!�����e�QB6g�BƲ $���_���+�8��ěY���e�vBA�4��+�NU�~��>�7k�LC}]���+�ѹLg��D��]�B�ӧ�\�s���[WW#ۢz-�l�%���
l	0��9�h���Ō��,�-�}a���e�¦fh�@����� l���^�ݢٟ�x8o�+��8�c�h����6Hq�G���{ ���g�5.$c��
=��X@c����3/�CΗ'���x�KtP�}{�<q���sk@���+���;Gtj|{EW]��r��[�������S;3�����}�6>I'$5�yT#S*I5$!T�_W:s�~�h3��
���"}�c҇�c�`��@5A�x+`?f�� /d�����H[�$Ƙ��?���z��"u�\u��fG����z�0����^����[&6���ab���7����<�(n�­ fC$.�LV%�w�:�zK"ʉb��0���IlwvĐ1�lM��F=��/��n�5c�.j���J���/��Yg\���&�5esy͞}�f�<0� �誨�Y�A��O6O���dw�w������k6N�b@J�S��H����i��h(�m�=�Ѽ�F����1� ��?��\�F�UG:/0D� �\m���p���w�AR���zb� p8A��G�M���#��Kw��ԳO讯.��\����L�r���e��k�~=��M�fg5�L
�*��Z��ve�lEO@�m��$-;"��q���n��"�	P�Ff�;l� 6�,R�LҐ��W��8��s#§n߃AMy8����1jGd��o\;�y�1qՊœ���j�Զ�zӛ�ӌ�����Jk_X�r9�c9E�Av�項���a��A�X*�j���b���ISC���$@���Q:3l�-�}��/+xb����j���V�.�L����׺��7��?��9���֯���mV��JnA�O>}�	'y�c�3u&���m�c �Cf�q��,4^�Ќ�6�k�׋v�o`6 ���e8��6�n_ړ�e:�$n}R?$�?cc7b��È!+Μ ~K|���`x '!�+@���6{�{��\�Y�?��p�b�̛0 �}�7�K!=��?[��.}*d'�<R̕t�U��ig�Z���T&�$�V�Xޡ	wUOO]�zN
e��jToY�<��x�7�����S"�����~7l%����L�!�a� T���K�"o��%�>1n�'�
,�X@�@��6n����������������ï������J=���1�L��M�Wo|�B��}B��	%g`mM��v\ǹx(�! ����ʧ+b�Z�LB
�\rIP0@څQ�Id��0�aet\��*�'z:~����R�Ӓ%���)�L��j�S���YU�7�����%G�$ LLx?e2ĞQ�х#b�f�]f�˓� ��.��l3�� �H��u�&�A������4 z�Gz�pߧ�f�N�73��P᝭iG����{b�3��x���a~3����N����u;���E&�8�Cx�� ��P�Dr��)����D���۾"��j�Kg�~��p�~�zT�R��MM�SU-OЄ	����������JT-l
���-s٘apDGX�!�@H��0^��g�&j�xӘ� ;��;����P�u#֙t+ި搩A���	<�ZO�����|.��k\;� �M��řkon)fX�ʔ� �qo=F�gLӒg��s�%q&�h,�`�B�3������2�ʈp�^\CHdF�
z��w�+��Au5,��7�blN%��`N��$���l�G~��֬^���^57eB"�fM���mR8����O �IQ��ד�)UN�3c
pܯ��-����l�l�=q�y�-\1�؜��k�kE����������h͜<C��t��c������
g1�m���/\�3`d>8������8v�wZVl�^���m?�c�2���z5iG���u\U�q���	z�Q'��}�s�������|�/�-�jo���W�#�X|���h����îC�+��G?�YT��a0���q��
u���i!��~�7 �aT���F.��Ƃ�_&<y��w6uo<&�Ԅ�i��l��O�*��]�b�։N؂��C[r�e,
�c(B'��vĖ�g��F ��=B5�5k��G���␄]A��1c�|*K��/�鬫Q�(�k���Y�WooWOR�2�d
�,��Ve0����&��هc��,��@y��o�'^��A(aČΟ{1y�/�,;������K �1�JV L�P����F `�O?�ϙ;��Pf�\k���/f[3�	��e�t�w�^Ω�H!��IA��6�z-��	���λ*_�T�q!Lx/��7��$Ԓ,&����|N��?��C���� C�ϟ���7�8���>��]���ο�R&cY����Nj ��󦒚��s�V�5�-_4���V,n���/d3l[v=�Z������POx��v�c>N���q,��1+�)����)1+����b���w�3�����Rc*y��6�%`pI�q�%��%1SE0��>�J?uA����
;x
M�/T	���Y��e4w�;4m�tr�Qݛ�~c�d�n]ş��nc���$�g�y"�8�~����������@<;�=5��F �����t��t{�S��g2\�m�G���� �t�R�v�"���.���p�Q���zN�B�z��!U���M���ڦJ��l�d�0�6'ٛ��x�,!�]���*��n;��a�=~0��y�w�DMa����xC�C����O�&^a�\�r �X�`�+�m� �dGP�'��ic�z�
Y�f���Î�34����+j! ӫ�\� (���z��ư30l� ��F�\�s���t��H�Â��f��_�������~WϯZ�lnɅ�Z�z�	�k��+��g4m�~*d�����3�<)=����%���qB[e�E�i�,��ʭ���{��i�|����x-ē��[k{w|�%�7Vc���U�v��QS�ګ�v,h�m�T������є)��cުw�C==���A�b����?��N��$d���u��s�v
X�6`^�3`6[�lp2��,�9�����kh�: l��^t�=�1u�w6uw�*jo�7z��ʚ2e�`]���mÎ	z�#P�2�Kl�;Wb��5a�7qa �;e��c��x1�v��n���r�AZY9c�^ߠb�������.��j�z������h��5��B���@8�����[2	�p�7�xW����t�3��dY���n��|�pO�������:	�^�	Cz!6}M����Gb�[�җ�
����������ޖ�{�{�f�~��>1C8Y�V�m4�IjK�I�ĳ�����m�x��/,@�M+�i�r��y�� ˜!��6b���g�p��3�#�Q<_�y6�\6��k�9މ������"�1?Y� ���yD���~Rq�"��gB5��`9X��2�@30�
O�1+-�5`L�^��B��Ya�X�W�z`�@�X(א��A�q��j��B�G--%m�C�
�%��_Tk�=�h�N�w��:��6� a�{���-�� ;�)F|n��q`/��13Jjz1�qrRr,� ?�	���o��1��� �e���L�8���[ߺ��4�|�Y}�+�%�|����/t�;NPw����W�>A�W�k�z��q�_X8�r��y�>��Ǝ9�c��U �f���F�����-��]�q�٤Ћn�1�@��;�I&;�:xŏ�׸�QL|��u�]7�g̑�6>"��5)[&h� �!}lZ(��8o��6Q�v�*fet� �n�]�C�>f̎�2�����ư�gN�I�A�����ߣ�v��c�?D�'��W��%%�q����*��� �p�ys�־�NW~+@��:�	����)1hDS~����7�12�j�1&�+��gZ���u�1�t����X&���Z��}�/�V*�������9��R�K�B�~��r���g5c�#��v{�^o��J�.��pZ)j<&�s&f�7h��Ldg�6�ۺm�p?P��8��Ƅ���B62��z0���]����F�]w�y? �㫥#�1;&Wj�c�=��8�<V�8��t&[*���3��}�N*O�6���1U�����S�A�v 뵒�}��Q_�����t�E�PlҳOm�ɧ�'��Y��Xb�[�^���:{[��e���Id���v_L3�X�̴=F���Gh����J��h�����C��بZO�γ��T�q���;��Wb���K�<���z���;5eJN�~�l�r�q*�K�����>v��Փ�G?z�f�<T�2R� 5�pO� �d�v����������Ƅ�ޞ�c5�r�5evmF�8�1�އÞ��S�����n�a���O�x~q{�/�0g���#��bU=9,�Vāp�q+F�:;ǒ� �w�xq΂��f oK���ټ�L�85 ��1~���V�ʽ������k��L�?|�cz�k_��˻4��w��/�Z8�4�rν�[.~iFb�ܰ1����w�(��!��x�c`��bO����Г�x��	$6��+1����Oa�e����x^��X�����4����X�z�]��٧���ޣ���v�5i��iμ��S�u�~B?���i��]4���{����2A��^g�_�<,5�qK�����):�T33]�nM@Lr�W/��egP������+^5��>�ûW�/��2��|�n���X�%sj���x���'�yaq[����ld�����+�����]c�Ke`J�Y��mS��O+v4������|f�EV�~q�>��k�裿R�(}��u��k��>���3T�4��9r��	N�7ڼ�5�@��̀��`�El�����ld����D����X��(9��]CV��Ɔ�-v�F!fk���EX?ӆ#V�4��;^��3#{Kq�ʆ����3���I��x��A�Y�����8�kƽ���i_3;��`{,c���X���G��sZ�d���vU�]�0��_v�N�}�:6v���\���
m��>��ŗ�W��-iܸ� �l�pQw�0;x��զ�U���Fh�~m���Id�\{%�����#BRvt�m�.�4�7wЇ��wY�Vΐ ��|����{��K^�G�_{﻽��Wk���ԓ���i���R? \�	�dan3JY����q�B�Vi��̛,T���꘻��1���d�=��1�1�z�!FݴR�3��Y|<��p���%6i#3��6ǋ7i���5����-�L�c�g�n����ux��������Põ'f���G[z����%��J����t���ּ�NPWW�>��O�ޯ=��^���ϿR{�}@8���4N� $AMn�W��u���A�����i����:�����%�S��M���'��^:�o8�jaœ4�vK���{�b���S̄c dW�po�.��|��kt�st��ǫPl����Yg_���A�>m&<��s� 3A�v�?n3���bOz����eo�@i���ǆi�g 6%��@�`�4;����wm,�GiZ/�&����u�q��:.���ٰ�š����H��c���4�r׻<"m�Y����f�Eǲ�Y��ѭ�W#ݗ�OCK�-��E�T�/������Ь�oP>W��zH���۵�#��|讀1�p�Q�?���4��$���s��z�`�n$|����0�Ɵ�=��0؀f���&��f��N�'�[��:9�Տ;�g�Q�qU�+aO������~��ϴ��4󀝕-t�l�������Q�:Y��,���ԱH���1� �l>�<.�9�k�� b��y���n=��o�(bvf٥�ᦔ5f�1�ĉ��i��������b&2T;�No�u��Y�~Y�}y="�$�%RiO��c٧��,6�d�I�e������D��!3����1��Z�sҞdl��bj[<��� �|ų����]Մ�y]qջ��YGhܸ�J��V���������M���z{)yYT6_V�ZQ��2�$�K_�� � l����H�X�{�P���5��_�翢 ���r��ń�pD�CVʴ0��ck���1����Daa��V�� \��Զ۶i�]�iC�RU���6^O=�^�x�ձ����/�0�-��>�p��@L|( 5Xx"yU��{贗X>�Ryp���'!���s��k�a?s�v��4��[����e���������:o����>�}�����C�q�؀�k�f�#M����^����Z>������>���Ǜ�x�J���,3��3����� �ٚ��x6�`�Y����>��$E-_(�T�	�w���=ڰ��9Wrr�1���#Y)S+)��6�H�9ֵ�H�H���M��Ga6kLY�zq[����@��t�l�(�$i �d�=#	j���<610��M�tJ�����U���d��Śr�>���[�yd�>��E�x�z��ԏhd5w��6mor��c��L�>�x�P�|S���p���"fαu
�Gb��.i���ń3��3hx �gg`����(1�1�4����)�!p��2`{\b6��}p8Ǚ9��a�5�vJ�A�v �Ά�����:�a挌Y�w���<֩��7��/�W��'�I΅���4i�8͝������Z�̙J�) oK�d��m�f�LQS���J���`��{ｃ�ͦ͞�B�)�wsI�����ޡ�<_w�u�t�Acw�\r�|z��FCeGp�=B�W���c�.���IY<!͔�(����Rw������a�������h�굡�i>WRSsQM-mZ�zcP�z��l]n�5wΙ�6}/re)�	dN_E-f/���7{��pb���}��J3]?�{CM�l}�(i��B�H(Ļ�x�����c���H�����H�7���oo5EnT�Q�:v7�vV���En0v ���N)C�.��i��R@�<Q��=���cEǸ�]����x`���Q����Cޜ�g\�ߴ��
��g�����/*��e�i����	7�b��PO���,5*�8��bSC��^�s�j�U-��:�����k�T���G��H�.��L(?��J���P�O�k��M�{S >�}t�s��B���	Xx�x���E����\6�"@t    IDAT �< .9�03-����SY�z��.yF]��SsSC}}��+W4q�d��Sn���
R�0�����~e�y L��2��� �!�%Č(�$b�|c@
h,���D�aƘ]��9f�~����� "��ras���K��ٟ�/n k�a!ŏ����8�m��|츞�r?p@���� %bx�Ϻݱ��?:D�U =�x�ϊNS��
8s���T���=��C������9I�q�Ɗ���U��<����̌�p��b8oh,w�g% �U�G�r_+��^ݠ��L�I[��TTSk���k5QV��ZhVo/ۍ��q�^�t8�ۃ1>>�}86����M��?��I�qɺ����@8��|���ߘ2a��<��([��B�0���I9A��A�cX
�,�5NQ<��}�׊D�< L^��{�A0����MM	&ŭb���[�1P��(�ٷީ���ڸ�O�Ţ
�R-�\�k\���ԝN��>���S�<R=a�>���A���4x[�.��Z�(iV�sm �ﲑ�Ԅ�a�Y�}1���s�x> F�*��� |�nP��ǹ_���:����� � ���\Y�y�S-p�sJR ���͐�5�w��FJa*ڈs�1l�g��ϸ����������h���Av(�� ������ (T�s"0流��G���m=�n��A3=��3!E����^eգr��9�/kVo_C��O�{�|s�j���M}�l�h�:�3#����/�)�<m���m`��L�^`���p�=2�Tb�|"	��=�^'��z��#�q���4PO���^{�؂���~h�Wߙ�XHKk�jՆ��ݣF��LN�����S�冝�1�E-BA��ꔫ�4%��A�if�Ii��I���B��̘1#��b ����G�v��@>_U�����[]{B�x�����>Y�>�<��7�I9�F1	GL�'�!&A�ˑ@0�2������l �FG�A)��Åtb�3[��5�$	�1�iv�{�:�|���L$�0��z�{ܟx�ĕ������R|�S�gr�����< 퀅`L0t�{�Q��Xo����C��<z	�@��u�6�S ��)�އz(lЁ���^@Ma�C�e��w�>���;E���.^�zU�����Q��K;m?NMM5��!&\�6i��u��ў�LW�RV�*e�.Ԝ
�$�P�` t/��2��#��b�9c@�c\���!��˸!_��(Rp=0�3���f�:��y�K�w#�����W_}��u��#�Lza٢���C�[���+�3�X����*j{�fO|�!m���Aa�f`e�H�d��Ը�>��;�4����5��E8������B���/|!���$�bya�@d��Z@�)_R��1�1ǙX�b5��<��]r�U��ͪJ��=X�=�1����ܟ� \��u�Pc����,���3��k��r�,>��y�G��	3�6�����0^�������� ,�8��(������\�������N1�0
�t�	0ia�0�ab9��w0�i���|Ǆg�>����y>���  @9 ���+���Q�T^�I��6��x �@tC»!����4�q�Y���[�C��p��O=�{�v�*}M�Ь�Ν�N<R���pe.ӦR�E����o_(��VON�A/���`��?��3/��<)g��7�9��c]5/��60Y�������1cl�27T=a��������{ǫ���l@���\sͅc
�3ϻt��/�\4�^9�R-)�ɫ�WSKKs �=�z��>������lM��lN�q>�7��(��Q� 1
- JO=arsY�Eh��T����[B�O������}3��,ۮ���T�8�+���o���M����i���R�@��Cج1�lM�w?�s0��A�ﵑ`���i �;� f��p^��ű������8��V�,�@76ʐ��bHc��Hߨhq��k]q���' $��K��γ�O�-z�'N��st�I�u���Ћ@��v�Oȋv�=��a��-�����29ai > ��_�@�0l�5,��q0��C���v���^r���0
��c�6Ң�Xo���z���s�"u��P{kNW]�>�=��z±�-�m��ڲ�{Z��YW&۬j� :l��K��.�{���M7�<��|�;�O<��`h���y��o�G���u�܏9�0n�/޸��r5�r<�x������"G�����n�馋��o��["�M֎ ��ٰzQ[����R���&���N����4Y�Oy���v=��s���,9�f}�a���Ą�pf��~����N�q,��p�
��<(?J}�y�k�UB�?�Ov,k�<x��y�Vؘ�e35U�6��?���ݮIo��Mݶ5���S�:�̋�ݕS�)�� ��i���*�bx1����
�X�Ǳ\�t�i��q
�9�Q^�H�2R8"�	�����@p&Ɵ~�)����7s�<��\ȡxU +z���5��	��q�y}���C(��`�.��;B��"��<���c��0�	`��:>G/��LpXυu����0fX/s���,��9j<��Ah�?!�{ˑ���� �乧�h�������Iͺ��s��YG����J����f�~q�㚶�Q�i��jd
�د����F������#dƸ^q���Qo�8�s�!��NcG� ���z��y�������8��$���{�a;�������Qq�8 ���~��7`LAxƅ�Mya�����'\)�B)���6���t��o�#�TO>�t��^f�h�]U��R� E�����s0��8��f�p.'fP�߼����x?����)[�8~�������Ї�SO�
�9�x}��sU(4�G�i�T)����0y��%������B�����p��V�����E0*�a�L���c�~�A�r�ӻ�Frg��c�n&LȀ��SB7ƞ� K�i�f�q̍�1	a,��3 {�9��yc ��|H� ����[�c��41���]E���B?�D�k�m������� x'c�w��ť��0n�H���n�ﳑz% vs��x>=��i�s�W��թ�m� �s��Je�~���u��Q�:Q��M:����y@�Y�������R�$��	��� )tQQ:� R�@B�Q�qG�QGfH�
�{g�5�;cEE�����S�~�o��9��rJN`֝�u���[���{?�����u����!G%�R��e���S��e�]�!8�b�40S�Pa���I�A��ڬ�3p}m����@�/�'�6�ߋ���q�8+�J9��>z�=�\7� <nժǫt,��nڬ�u-:����w�Y��z����ٙl�G͆��X�3o�#$�iӂ`~����b
6�Z�`��0ر�! ��1U𽽬�ۢ0p���U)���5���1=����k�F}�>�IS�虧������0�#*�L��-i��Q�'�[e�=�A���o@�
m0�s��km��@�s�n���¶����{2pa~ L�Ś�0��L �Qz}�*�E?-'�況P�3A�����Y�q�#��JPl��͎K<9ޡS.�ͽm��;~g��Y�@p/ƻ��k:r�c���B6��g�s�"��+���e ̭�������K�葇����ujn,k���u�Egk��պ��껏=���?X�}t��r�r� ?t	iJb�y�<�@_��W��6p�g١���?2¼ cb@���l����y7���#ք�X��i����X�ڛc�{�k9�N�:u���Y�|̠������?�е�X���">�g�q���6U?��h���P��0����a8��cDg�Y�`2��.x���E0<�C�0@�{X�:���zo��jG`��li���;tӍ�ʕ������go�[�v������U�U������9������Y7xt�A1��	���OWA��L�׈A86G����x�̭��`7Р�	�g�s,� 6MLV��@�Ƶ�m~q�P�ν���ڒ�	/�q&��;6�p?�1cԑ���dd3�ׄ����9���Q�C/�\�~9���v	 �N{��X��皱���s+C-�C��+��+_�??�U�^���h�7|Pg���ڸ~�n�y�~�����u��kn�aG�R�$�K-�F%�s�r����!?daYǋ-���6;X</��wh�<�gd�Yg�ٓE�9���>Y��+��3���g��= �i���	L8��<r��wlXA���u+LLW���� ��艺����Ц���7!D�d���6?X@�$ L��A�N��P�PW��>еM�	�c;jB���>X��dprj*��#�*��<h��C��RG��ϿI�-�������Kws��v�<�
��Qԝ���t��P%j{KY���0�OD&p���A�,�����bu���|��!е��&llN1��J��6�x������`WM
$9����`���C�T��Y��ǹ����E���W�C�`��_	g�K�����s�Ǝ�n�s�{���U��/�;���Ə?P��Z���jsg���Ň��(���15<���}�� �L/�>�&*k���b�.����p���P��oN��^`?��o`�&���D�Y.�[�VK�l��;��������l�w&:b�����sgiźez�O�14 t\�դ�	 �ax���N
�;2o̚=�	%���k�q���� fT�/���V��t��1gGV�a�WJ*tm֜[?�be��=�T}��3B&Вڃc� ��l����9"��3��cbS��3���O
��|��a`��8���06ؔW�X�1P6Ma�m��?@4`1��ǚi��_��@����w�cb��5�Ʀ����#��tQ��;��+�e�Wj��_W�k��[*�w���5�=*:���	����В%4�_k�}�W.�U��{�|�a��::��
���%�\4.�M�Ih�?��OA1`� D�s�	6\L���ڷA�"䎨�X3�0�e,d����R.���]w�qð��W�t��+��7Wߐs's�N;�T=���kɲ�!l��au�����@��`�ǃ@ '�pBx(؃Kj�4;c�Z=��c����q�Οv�i��.��%�os���-���ҟ�����cu�Q����|OIK_�Ѭs�VG���%�)͜y~a�\���µ c 4����w��?1Ǫ��A�ks/<Vsm�����LX���ju�{8���; �m��N�Ys/�^�G�5���s{�����ׂ�`�>>vG��ζ��8��h�zh��
ɦ�7�tipp74���Ӛ��z�wK��>G��q��ne�Ⱥ���T)�T*&Yq؄!bk^x�L!bD�xnجd�/�;�gy�[���0W��=�v�����0�
3' �{�89�lF���6�';1W��b6���Mw�����&L�ܸ�5��[�'c�舷�&�z������֮_�j�B�b	:wG��xP�^1G�[�����(���
��*��w�}a�
D���g�\/o�9"�x"�S%�/k:M���&˛5z�D���M������`�% L=a2��L��]�]���� �An�!FFqh�@��L��l��M��`�Vk�����^`��MO��$f�Cɥ�����5�m�����p?�9�K�J�ٶ]y���z�٧þp�Bݕ�s���Y�P���U�~��ܬ���^�ƾ.��\����A!�����&-��5���D��BRc��m�D�x<:[��v�����2�L ��	���1�W,���}cre�nظ��rJ��o�}��ӦM�8�P;b�K���g����<��t��g�W��^Z�2�1ǖ���A���#�!�=8Z�.���Y���r�uׅ����}�J��(�m���/�� ��@�-�m_�p�Gi��mzy���Ve2y54)0��Ͼ����_�ё؂�a�C'k���>fr��D� ������13u��P�C�p��X5�Y�ꟁq��
���MW����Ү��L*;bnٕm|-�m^�jY�Z*t��Tt�������fHDO�(��yO55�r�.)ϙ��A!���=}�����`�2����n"�K�1cF0;����{��̙�����:����;�@-��B�YͿy^r<� �p9��磏>����t���΄]E���9��դ5���4s����y=�̟Ö�v��c�p��!AN�Dh��@�`��}p���#,�3+S�Y�3��6�$��1 �U�]:SQ�5������6mH���*��qcv�K/��Z��v3��؄��>s�4�J�ⳳ�~zU��E���t�9��[˫?�i��sG 8�����֪ݖG-�0��YR�:_&�� �Kj��4�������l��*vwh���ҩN)UPW���B��1z�)gj̘�T�Шb1�J)q�Y�1�ݖ�3���μ�|@dy����GG�ܘC�B2'a�c5q �դ��O�+r>�&�{�������.��JB��j���w]���V�؄x�~:��)�(����R��x���6���z�bV���P�6G�9���{:Kܟc�<�b/?̖�!(�:�q��*�h�吨x2yңN��CJj9�wu�I�L�:�Ⱦk�a"��:w�y�<���A �)q�ݸw���1�:��H��;�m~qm�y��1���w��A#��Im;�N�u0������<�%��xQL���j,���ᯠ���W.��a�L�	���\���TW?N�BZ4I�'�|1qd��5&s��^s��z��fln�{�Ø�$1K� ���;���!a�1А�B}��_��0V1� -����&#'�6�J'�!j�̷�c�Ǐ<��u;����-���=E�6jB�	�a���o~��M��c@@x8� ?�,�4�,��:�<~#�{�w��� ���Q3D�I	�A��2��y��8�!���,:�&��B�[�<��
��rlwTج�&���kR���p5�J*���,��w��D���88� b��<f��q�c/���1�m/H�2P˯���}����<����As!��ׄ�ϵ��U�Ȅ������3=�yf�����`���x��C�U�$@K��|!�l�I�N��Ɔ&�����T	W��E�x,|mj8I֠��F�4,�^��l3Z���`8�v���a�0a��!m�9���F��m�Z8!�d��l.�J�\6��=��9���W���4�	7�7��Q�q��3��G+^Z�%/,U{{bǵJl�<�l5��WNm�{-�f5C����k�C���W_�C9��%��	� ݡ-�U���1�[l��Bq�~�����I��Sg��~C�ʩ�ҙ\���3�Sʒ*jea�I����L��sF$�jI��dj�X�g�v��;锖�\�i=���w�j��G+�KJS��U�u�m�}u�1o�GLS{GQ�JJ)�WJ��i��������R��K/�4�p�l�/�	��~!H�9��)���p�{�w(h���66�Ӭ�cC&t�����ߞ;w�u��c��qkV?4���V*�:d�)�������8I�M���Ͻ�ի��q �M ����0`�}̪��V�">���������b��
�*F!l4_��8;�͌�cε���*}:C���*�4zt�Ң�h�2���x���o�jU��� ���0�r��3�Wk��gD�!�W
�.Z�@ULu]~��q�)j�˨��H�Ѫ���^Q*3Fi�V��R%ӭ\:6�����Ct��E4�B�3gN��w�D�>�8߉~ ��sX  c�.�1_��`Ä��DJ���t��Cr�Y2f�6>B    IDAT&��];Y���R��调�����	Kt;k���!��}g���l�֭��}6^Yl�WV= ����P������v�|�PҎ)�1o޼p�PGTH{��߮�|�3!J"V�$f�-Ղ���L���l�F�ɨ��U��l&=��պ䒏�u;4�
��JF�g��)��1W�R�`����pL��k�H`WH����5�������h�u=�3�ÚuJA�,�њ�Z��G�R�Z�^�|-2�����K�Z�,;����>��`������ʃ=���������!`�kӣ͛�/����Ô�(�
^8�ӱ���W 8x��_�"�@�l`�Zeg�]»mX�P�uô�� 8i��V�iJ�I���ScƌN2�÷s���8�֋3&U{,3�_�g�(�DG �ޙ��B��te�`����C�j����L�ݖ7nX�_��:���:��7)�Mj��y�K���Zs��E�% ��1�P�	�����
d��&�W
����}�+�fRjn,覛/���:Y�9�TI뷿y^�<�J|�&N<P�JS�쳱�.D�
�`I�� # �@|�C�8̊��d�'����)TX�.	 g�9��q��sc �?������kሃ0�&*�Q�;�7�R�T`Ι3��ag�ׯ[Tױ��Α��-�C=�jW(�<��#t�'�% H�H-�l���#�P�����s�y�sQ#0�� ���:��x�� a��Pq@s�6��� �J��u�LݫB��>K�&�Ջ���}g~@�B�*���� 3f^��p�3�g�`^�WmF��hD;(�W
�+V,�c�������-��NU:UԿ������Y�^���O��1ǿ9�
W*�����F�f��0�ǹ;b��Թs熞�9����.�x����M� �DcqVᓊ��#ށ����)�@���E��.�qkW/_-�@�#BԚ٪VTH��DB�:��nq��,�S�(BA�t���PT��8�թ�t��2樂d�`�5]@���  �`&�ӏ���s6��hR�ahwΟ�g���&�у��}��[�?�R]xUH֠�O(����3߯)S�Y�M��F@xg����m$�J@���M�ڵ�ScG�t���k��wjs�z͞s�~�K�P��n��Nt�a�(�\}���d��#�a�c��Z�X���wp�S$����q�|r�q0���D(>;m[1����ua��;�Zda��*�e��4�8[N�ӏ͝;��ag�J�
�`��$麥LA��u���ӓlX�-gX�xKE`�-� /�W�w ��~��E�Q�ױz@�v�@¶'ՕԸ�w�������	g��ޭٷܨ^���������c�ЦMy����U.7�,*>�͜y��L9<DRT*���8i��H��p�@��RwG^������Ӧi�����Mw�W��V��s���a�&M>\)j:gɈM���٤�3�"E�Al64��.�|��7�u���8��q�`��7{�p�5Ny�k<�b�`Q����WųV�Ȱt:��.��7�[�n�xbsKc`��1WW�Ls�8��)D@.�B����u��Q�K:㒌��p�w�:�Շ��pC�\[4Ǻ+��&��j�^&�V9ߣٷ^��a��^���M:�Ѓ�l��:��K��7&�,��`��9+1G���4��3S��.x� ����z���RW;󮬹�]��3OQ�{���>}sѯ��}&��+����NRO1��!	_���͈�\a�q���\O��;v��������l��̆�̵��qDD���Ys<��,�h�kJD �zX�����V.j)t��ڹ���	��	������$����N���d������w�WBg��0O�	���3��.�|����k5��k��tj�y�ꃗ����F=��5��k��ѨR�Q)�Bh͌Y�4y2;�ĖOU4�W�17��C�8֫���7*����.��9fq�
�0��5TD�p��p�^�&Z��uX��q�'Em��c�]��>�~��,�=m����N����R�O���~���};�;`�y���qV����{�BZ�u[MB�w��0��'�Sr�!r��Mrh�N[7PL8�6����΂0��d�Z�`�J��ru]�u��������e=����_��^x�U�l��v���^�^9�;���/�����1i��L-���1N5�|l�O�����׋�.Z�ݖ������]�vQK���0��qN����������5�<p��W2l>0aq�m�����3��!��I����qi��vh��]�������Q�JS(>M�f̚��p�'��T+u���A�=q��n�\�Zu)��S��"��p��<�'iF�G�h�������l�LV�8�k�-�1=��Xc��xΈ��#���/0n?�f�p�'�.��@j������g��}�N���~�M�+m����<�6�ݬ*ŋ���ŋB�:�+Axي%!v�T(i�>y�L�q扪���֤��m֓O���_����J�:��C!����I����W��W��ߛT��oG@ئQ����\y��NL,�g��wo���+�u����X��'Z �>�@q�H��^f�NQ68 L��	q��y˽0it����=V�2��mVS�h-{�]g�y���f�������A��)+�)�*L���꓋ۛ�=F�q��/���;9�s=x���:��LĬ$vV8����w��^f���t𻁆�9�����r?��+m�6��?�q^L�P�=Z�4�\����̺�6G���g�jp��o�1�������Ƞͽ}_��>�{�c݋���0ǹ��e����scW��eID���.�4K��r�f��N54�U*d��쮍Kjo/�P��u!A#��͙�b���W��7_���gm<������ZY� cW̼��S�����+�9�U��|�Ec��'_��v_�jѨB�I1a�[8�zŝ��TK���|_���\fC��9�7��p|ߪz��vi�j�H�bSV�j^�BU+���K�/����*U3J��	�8W���5�����d��3�����d�i��'�A����,��!+&���kX����f��z�5�̽�Um���l��p��f}6�����m4�Ƌ���'&��^n69X}�/N����	䁺o3��������`��˱6�Y�f��a�bD�bY[�q����V�I�A�>�Mܖ�����#���bL�Au�4~L�.��]z�U�E�D�R��S}ݨ��y}]������f�&c�d,Jxq��3��qw�ׂv-��u��{o[�?��+vc�Hᜪ�	ׂp̸̰�[���9H�����ʃ�5h��vA ٢�c�~���Ժ5k(�r��r�z�*�S�ohQ)UV*]PEe�
�#�-���(��ʹ�K�<�'񍞔V�a� �����4�&����ӓ�L$��a�-j5׌ˏ��!k�~�y��<d0λ7��b�N�`�um�6�Ӷt����ك\�u���݋�˪���=��1+�6��5G�HUl��d��W;��3}����!O|�u1]��y�~�����k^di�Uk�(l��UL~�?��GWV-�hۨt�]�P;K�6n���{�Oz�v�c/e�.�N��t�Du�)�6���M��˹�������cR�������~@��y�Wu�Q/�H[���c�K[
�0�~A�6�n,>��b���U�xL��~haN�r����sO������IM���F�lV�RU��8�U@�"M����[� ��;k��h3��K�l��$�0Q)��>1	*�!A�	j(a7Ȉ8I�'��_(t�9 $��Z�����'� �qA���d�=U�l��b�]p�N��dbq0x�:��ɉ�Ǝ?ˀ�L~��K6��L{�;X�Z��j=�|Iq �+�^C��I�B;�XDlF�:�[& Km�h�F�i��XB&�.���m�t��yCO��g �\YA&X$y�ĭ"/�̟Y6ϖg��[�ߕ LQ��}�U�lST%^2!r�v��봹�K�:Y�l�r�d�qU*�{���	O��Z��s�x����rCͧ�߇2G��%[1h���]½���΂��
k üϷ����b��̭?&�C%�7[/�淿P��LU�Rw�l�ʤ���5&@�) <�d��a&7���%�� �~3��8��p���0)@��JR 79�8a|��\yw�1�9 ��K� �g�@1񩻊�)�xҖ_���xF�-���m���B �v�`��I��Oo[*Ϙ
ZLt�B�8��}�%�˽�~�\3��~�0� ����CF�G[��"O�I�*�����!��ܗPo��bĽ� M���:,X,T���; ̋E���vȀ?τk"K@��Bv$, /G}�4�+Ax��������J^jl�W�ܦ��M�$ �󅂪鴎<��e��ZM�.���WM5�.y�8d\ׂ�@�n{�����������= <��ˇ�9�Q�)&<��QadC��b����1� �؛��\�kS�j��?�C֭U�ܥ|E�[�M�ղe��kV����J �`���c�2Ø(v%� l�	 ;X�?�,3�aF|���9�&�yp<���
�	l  P� HS^�: nP@���H6��`��I�
�'���Yک���Ϲ ��u�v��~��<ٶy �̖{q-&�h3��Q�q�S�C�],, ��� <��*,<��s/��>Բ939�Ŏ�xN�'σg�,���^ 8l�c i�N_YHXmd�,���`[6�;���b��<{�gjA��^�M����c�}G�.JS�5����&�^T�浹s��~��z�[߭}�>T��U��3���9v�B��l���V���s{M��.B55��Z3���]f&Nx��+5�;O��φd�TgC&$k�����r���<B1(���*n��U:۴�X�G��"����L$۸��Ô��;?<��L�#�>w�)�U���ՓߨƦ������*��Z������Y��z0G�5�bM:�e2d�kA��2�`c�!�~� �l�]�:1��<��L~ؔ��Ӏ�1��<X[G��#�r<�@�8����y����� X�B#{���\� �xN��H�7���q.ㄾ��{����?m`���������S�9`gq��� +�8�|0K(�A.Ț�T�b���A���� �bd�����>g���g��u�xq��;��MH ?�ݶS�a!`Npm�X�I�,c��{7�\�bqp�mZߪ�v��}�l���ǩ���r�G�ι1ڼ9�je���VWwYM�Yu�t�:�����Q���Qf�|�]܋��X,s�`<ύC�)��e����������No�����4�|Otļy����/���ܴza}��̦Hs}5����P���Jp��q��OT�J��{6�L
ob���*��t�Վ������d@�v����������	�Þs�r�z��Z��S]t������^
;̚	���Fv�M� l0 &�6��H>��C��N�(X-�������W�@� ��f���0���G����C��^`ŨͰQ��8R���X8�@���� �˱�����xؓ�aV�7�����X!;=c �9�1ǀ H�1o�BΜ���&���ڮ%���{ ��XlXt�&�&�"�<Y� T�@�]a�L��&���dK�i}@saQ�"_�c¶g�"���ۆx��$ WՒ�/�-Rg[�Ǝ�j�͗�BX�t�ڻ�4n���v�mzmr��Z���U�b�++��w[6C��k��2 �w �,���f���LМ�#憝��a�&*�D�d��D���`G��J%��'|հ�0{��~���ζ��)�TQ��O1�W]CN�<�+%*��� ��#<Ջ��g�B7�5x۩��v�#`;U�jq��"�@�d��!?y�3n�~���j��M�[�:M'��`Vk�t�S�	��JՆ�w���5�� L�"|wu5;��	�2�=� A����dE^  �= fnL| &� 7&7�s`��x��+0cB0�`�� ���po�wHh�L��6/ �q�[�\a�,V�9���l_f�� Ф/����-Σ=��x�^��π0� g�q]Tz��
� ʹ�``�˸����3y.��p��EF�l����2d� [�s.L��3��3�9�;r䙳��o��bf*}�0h�:Ni��%z��_S�R���Ҝ9�駟�;�T����	=��K:d�������Ss�u�t(WGQ�d�O����5s5˷&l<�fc6���M��/�\kb��	��$yZ�&��e�}�	1G��r%��~��{����-�w_�baK���lu"@�R)+�n���'L�-�؀R�H�B�L�o��V{��v��F�� �J8�Sb�39 ہc/*�������)�Թy�����6o^���G���7d��S����_����JҖq(�% <� er�����Ң � Z��3Fd�V@��
�,lK�X�C^PX2e�H��°sO3E �g �ƦG� 610�l�@��!6Q �k���}��2 3�M�8�>9��`˽�D�%@� sM��Eơh��1���P��	�v���B;+���`��]@��J�3����"�2�9y�Ŏ6�Ok�Ȝ��\�5�d��	�̐?��5h� ���y^���?�+�l�KAx�KZ��UK�Jk��Ϳ\�{�z���ӟ�J�7��|OVW^s��8�DeӣT�H�2�T({03���GN��y�hO�ƳD�@V��ĵh<_�<�d��r��q<���D�geG'��:���W*�
Lx�A���n8d��Uǔ�Ǳ�Z!_
�,)��^h|��@M�vb�`GC�\<�a	�AD�a��n�4�z�:������78T�������N;P���f�m<n��ݺ������뀃���7�z���/�×~Lmm�p�Rզ^&|^ �lu
�}v~��&��ʢ�בpV�@�LP~�%�¶+d�JS�=�vu_�l��0��'��sڬ�c��)���ن�p��{  fl<&�:�~�xb0������ar�x�~ Q�f��G����1�Vo���N{i��/:|v�/�O{��H�s�#m������<g��$�����lwx�e�}�䲘�f�5�v����ыK�롅U,nV}]�����f�|�6ml�=wߧ�}�7�m�7�7ݮI�O�]=��R��d�Ą�{ĝv�i����(������a�4.>Ƹ����7� [s�Y�vf�c�@:x�g��&�q�K���{A��ٳgo)K@xb뺅�]m�3�\�	
y������+�q�����eU�����gM�`m04'��@C�`��j�đ�n���\F����g6��Y�A���C~%�|gE�n�E�?�+e�6����[O~��-[����a�{T��$LX͚u�&M:X�\W������=�j7�b�۔c�*�M0�����;	��������68��N�>������v73�Ë���+,3:O�x�q�l~�M��VK�����;'��teU���Y�q�9����30����m��2��W����Am �Z �Uf'����8b����8(�}6�N��6~w�`����#vx�c�˖�������o��	ҭ����N;I�m��9����T��{����M=�(�yerITQ�i�*j�02@���;�`*��8ϕ�Ȍ� ���������52��*�k��XC�q��@��,�D�`�w�5��s��t��a�Y㈫n:t�+d�[��A�!�uww��o�K���m����i���a(m�ST�Xږ��6ͣcѓ� � �O�l��7T9>�+_	v�3�8#�!��F������ǜ��+OG�    IDAT�+ ��ڭO}j���ԏ4i�x��wh����3O��%L���T�և*j��9��!�vN��.6G�m��N�X��@��6{d��r��"��;�œ��s�rA~�4l����s�����3�y&#���ʽ ,��g���|���Ά3�X��Ȃ����U_&�ߛM�U#{�9�?�JdO>�iƖ��N!�B�9����=�!��Ym�4r��zA�>������{YC�Y���SZ�b���Ejoۨ��Nͻ�]p�iڴa�>�/�_�ן�Ҳ����'t�qǆ"�
�d[#�Q�p�9��o���l�v�7�g��}.�5o��0v�����O�<L, ෾����*X���8��X���q�E8"�x���[���r&�}��9w��i�h�G�Z�`�JǱ�g�������t��S��w���Z&(����O���)�L�1���c�;�ٝY	��mo{[��~�{�9`G������������I�A�9��=�R��n�2�c��X�]v�>r�tuw�h��]p�uj�{[M�#f]lI$v�����Q�X�/��<t����'��fu� n���,/��|�sl*�y�A��s4��e�@����ф.d��	�1b0�������@;=�j�7�r���%���k�6��k��rl�����w�s����}N��5,��vm�#�ux�ŋ[��A:�%K^5���E�4�u�-�j�̓�M���_?�O��`�,��Oܦ�'��ik:$h�v�9���S5��1g:V�BB>>�<�����*����
��9�6f������9�@�߇gRL�e��t��;�뺩S�&����4m�L���������:{��Gu��}�;C��~��:;��
�xŬ�3 pf��`KF��>�h`��G��X_�@�%�53 �=�s-<�cV���chS�"���z�ձZ�<�kM:dM:l/��}�z������nVkkZ�*{�I���2:k�E�t(E�]E�]�� ���<�v>���F$�J ᪖�X����ʥ�V���C:�ijl��:�z��.=�41�j�}Qk[���L����جb>1���	���}����H,,���4l�̗���}�-� #�r���hD��W���	<6=،�Eڡh^^4@�4m|S�F'�(���J�J�\��;����
�؄'��]P��z<!j�i�6��N�!S������/�PHV�����%�ۅp<������?6�X��a' �����9�;Ǹ���5����إ����R�s����ܨr�S�GM�_�ިY��PwWV�j�7��f��v|��Z�gϬ��tF����.k��%z��QCz�T�М����oR]}^�tFݝK��W:�"�T�dT�P��v�b���0G`jt$��ؽ���`���7�	0��a��=*�^1{bv�s�5�X��и!�6E�u6h����������RK�l�����#�<rݎ�A�0 <�u͂����c��e�5�y�>��KTɕ�_��Ouw�H<��Vt�^fb���x1n�i�Y��P� gױ���TΪ��w�3���� #�4�#x��n˱3����nuu�V�ؖ�vR$k�U*JK�n�}�}]�6��	�>��532G`~�-�/T�1�����#Ǿ�0���/z����zM��%}����䓧�P���J���,��'�\Ɇ��L�M<��3qj�",�M{�ñ_�)�NҲ�Λ'{/��$�g��@�W��::�� q�|��l�	�����a&���OÄB���e�5o�m�s�1�w�Y	�c7�Z0��}<�ly����^�v�~�įU�%�/Q�a�?²��6A��*d����'}�8<�
v�����á�V'�Թ'������ Y�X��?�ca`Q�uVUPO~�~��k�3�UW�S6�l�Ġ��(�kR�C��I�U6�c;�R|;"x��@����;z��G$�+%`^��y-\�U�Mj۸I���'�|s���+956NдN�!�r%qВ�L)K�r�]3��π���K�%`i���Q4` ����7���XjL�\I�s�CS�l�4��\���8�,<�`|�;�	�'LX�\.�y�n�İ���+>y0��K=�I�8���u�Y�ӟ�{R/,Y6��� &:���!^]Tg� l������P; n:H��?:(������Fx\�$�jbo:�?Ɋ�.E=���*tC��J�;ܷГR:ۨR9�ԎH'�`�	;:"��� �����n���~WN��k�H`g$`~a�sZ�`�*��+$tmV�ԡ�F���PS���>5z|ؓ�2���$�48�z��8��sDQNl� N0�a�~�l'�v����û����\Nہ�>9d]:���o;|a���G`
\��.��A�j�C1��,�3��O+��<q͚���]Ӽ���'�E�z�;�ğ���V�8�L&�c_1�I�\���Kh���C�G��hv�qM �&ah�텈�`�#r�8�/��}�����"�=��p�t��?<�[{���,;T�kP�T�L�)ls��IBj�c.DG$�<Tt�P ;�<��ᶹbg&��9#ؕ�cn��e��N�K!���fحF��:��6�\M눩�(Wר�d߽�IB�P�$��[��Q�t�s��/��hѢ>��a^ޘ��8j₩�G@ؾ!;� r�����7�����IGP ��_Z�d���L�sn���7��M�g�w_�vas�sZ�H��ģ������Ǆ�e��T�0������E1�F�����>��!��f� 0�������#؏|�#�1�;�aV؎�f�i�P����@I�mՏ�oZ�f���;d����Z�d�2��O�	' |a(�CQ� �C8�2+�*�@LyWN��k�H`g$�5s˖�ᇿ�R�K�[�j｛�Ғ�w�[}C�
���<��������8V�=��	�h0G�Qi���cg��~O?��!��㏇�(�*k��8�YH�@(,�3;���9��	>0aGރ)�3�=��Ď�a�|���V������d�}���e�TQ������@xʁ�4s�=��Y=���}U�h(6a�ZbػR����Xe �L���0v!�;��L'�w5�Ky�)���i�Ɲ�e��1ʓ�̹q^TF+�6J�e2��K�K�����/��;�����*��E l��+��#������s^	��a�=�P��.ۭ+������ְMXH��ꐪSO���:5տN��(�kf�C�H�Z�`A o���>")�=d�X�D�M�x���;kҀ-�	�&�i!��%��q��tl
�0�����,�=��#jk߬2���.e�2߸��oVs�ԫ�?p��u���'x�Ͻ�碑.�0����~a.W�b���@��b�;��-dG*+a��=�	�� m�cUB(mm����Җ����%Y#횟}�R��Tvj���l�ޣT�Ki5���/��z��X	�V�	�9����\�{ߎ*j��)�0{�"�O��":��<�F��T�N��~5���=HF��e��B�j�G�M%͛w��>�uv�������+sZ��S��8U+cC��T��7"D-��>�����8I r�c@�;8�����N�ҹ�dġ����8���^1���3|��`@�&� �h.H!ף�z��.es�o�y���k� <f��Ec+�����!jg�}��;d=��ߪ��6��� �� �8V�^J��� ���@h�|�^P�9���w1j���"D����W��+ck\"*�#%,8�8��ؼR?����v�[�v�F�\�Z��[g��A�J�U�6&)�J' <�PeȘ�Q<c�ڀ�� a�;j}pL$���!x�}��#�-%08�Z�R_���*�ݡ���n�w�Σ�p����v���詧�뭚0� 廉��R�+��$Yc06�?~b��� + 's�'~v~,͊���7�9E�0����s�{z�?��ݗ�����	�v&&��`�����^?Tf
)'Y�;�nXA��5ƾ��|�	��LȘS?J�s���������z���a��}U�輙pl�v�\S����&8�!ܦ
۔O�&LX�� ��[�� �̜��Y`�0a�6�A8ؑTR.]��]�������f�#��
B�ٕ��>���T������i��I��5U	�4ү�����������Z�r�82A��#�	����/_JY�-Me͞�A͘�%�����|�a�ZӮ�o�SG���aB6��	c���K5 ���NlvJ��|���aV�h1?��o��0h�o��D��p{G��d�E�l�4a�9�{`��
6d�h�إ�z7	S;"��}���f_7u�Ø���ؽ}ݢ��'����F��رct�ߢ7|`��t���t�@���<w~c#ƏB� 1�%��x �f��}�C
�
��������?ݷ����4�v5���	��@�;���Oݡ�����ܻY_��{t��x�K������NtD�T��a��?t�z�����g�_Џ8�/�3���\t����xG bk�D�����t���K`0���׷���ݝ�R�-�߯3��6m�ܡy�>����/=������:h��*�K�P�.K텭���˂��5�*D�9~�m�з��H��Ox|�B�E�a�(�f��2�_�yET�\����a�r-k�f�0i���&RI�F�%[�Z���G��'��Z���~"L�8a�@���|ԡ:���	��+^�[��h��i>�����go�� 0�r��O�� $�>���"?8�"%� *@��j+�ج�.��,�RU��K��t��y�w;>�z೚z����3.V��S�ڒ�p�N3g\��SV6[��U*8�f��a(���vad�`r�~ ��ih���^Ԯt�.y�����70���Փ� ��Y}��o���U�ZJ�u�t�9����_�u�ݮ_����������?�9T�G���Nl�ٴ�����'l
��
iD*�O�_��onn�-���hB\a��m�Acv��_�4�'��wQ3��b��&,�u*~���e�ד�J]]��[o���iӦ��؄ǯ]M�Ɖ�	��a{�t�t����أ�Ӹq���p1�����?��`�&�a�AG1�s\�+k�1���3�LJYb��f�\�LV�/|�AE@�<Xo�Dz����(��on��j-_�gM�����7j���ֺu�:����z�e5�4��A�����c�)2��ׁ�6��4��]/���D_-�Woҍ�iD���F��|H����TԜy��Y�RG�f}�s���=�55�^�Ι�>$T#ĻB6]xU��}:0�ڍ>�1G=a���-���s�����:��#+�〯Am����C� ��]��%P���� s#đ�9�V>;�ӛ�Q����% <a��cʅ��ޜi�mη�yT��2U�7-��l����S8� V^�upN��f����F$k���7�G��T�{�VI��io�{1�ݖ�b�v�؄�֍��ݬ�z�N��מ��ԟV��SG{��j
�`�9+؄��\�u��N\�W�-R���"��1¶;8ݵ/���`y�H൓�� �l��zh�u�5fTJ��z�f�z�*�.��W�>���I���[u蔣�1M�1��d�^��0�
3�ܹsÜ_�j̀��������ĵ��i �d�;��8잏 ,ٿ /�؜	���L�0�g��qŕJ��9��[o�5Lx\�xb��
�d�D6�mN����1�����B�Pv�(�����xl2 0���#��@�]�B�	cv�m�qp��5�KF�6y`G��υ]<�쬑�1ݐ���_�{B���^G���:��m���s����؄{�VΜqn��H2�
�i+(��A�v�N�	�xG�D���+C���L#!j�4�Ϲ�PL�9-x�A廪7:�o�0�ՒVO��5�
��/��>��Ɩ�JSE��v��U%D-�Y�?f���p;s�p��͋`�
���?>�)��El� 7$�k��t��ǥ-}�XomD�wo���@8��>:w�܏�n�DG�ߴrQK��D�c�ʬZU�2�$[;1����!旕��sgX� \o(	Sv�84�������5RFWWO��^�u�{OOWXA�	'L;a���`�`�-w������Ru���K*�Z��6�;�*��4�PN+���sfhʔI��Q/�=�Q3�H��i*�8|��r/X�����Ȏ�F$��I�NHQY�V.	i�]my�4�u��W��oW:���fG������)��Q���Ja�V�$`�4����,X�Y�%m��k� 1��j���|M��/�7��p��zY�\�;��r��^����o��U�J���I5�;3�8�
��&Pώ����;4������ $�"na�ɞR�0��1���q�^޸B�\Y��V��W�I7h��n�}���^U�RU*KX]Uӧ�*���M���ԃ9���AB�9*����x�����H�l@y�5"��N�0�d����E��OiTSV^��t�a>aehl���T��Ln�R8�S9)ݓ��R��L�1�_ޜ��Wct��I�5�8�y�\�ak�6#�D%�b�͈��7YuXm|_��X�N�ӏ�~���+u����n�b�b�DG�Np��4�g�!W;��ǳw��ةeAqm����������?8��%������P��nP6EUa���F�Z�I�FOT�RV:���Q��;+=a4�8�@v�X�Y<�5�xa�ܯ�$���l	©���X�7*t��l����UU�Š92�w��u:餷j�}V�X�bU�$Ta�`g
"����-�y�0�dk4c��9�j��kƱ�����9��սE�|m�g۲ύ�V|=��L&��m��v�����k�*t�4Ä�ej�T�& 3e�h��r�7�c���ʎ-��8��1��Ât57/tX5SE)�YO?���=�P/���5�K���ZT�H%��Iv��sH[������PL�jmÎD��O~�`Ba��S�Qر�&(����#�m%08��li0!T�%5d�JU;���3� �f�l�0f�z�0�5�Tr|p�=sɅ����1�=c�͵ф�1H:2��ʿ�e��1q���s����L� �N��3����9�U;��M��|�'��}ͪE��0�#P'�
īIl����U��lA��@��<�=okU���!j0�r�]O=��
I��}�
9�ꛓ�wҝsd��8�����O+`LD^Yd��h�XW��f�#{��	��%˗�z�*���*aa�ʅ��Ad)�ޤ�R��@Ө�*���5%��{#h�	Ywwg�Y���f��&s	~$,�6_�q̌�ƌ>���p�&E�|��Zm>&�����;���W�)e���#���|��ի���X�A��qm���Z�N�	�(f۱m(�	W��ݪ����ڸ~�����rwO��+��P+�Q�J:ط���szm��Ʉ=` c��������Ӊ�F�v�,|�q�#��cF$0��&���p�C*vQĦS{���1Y�H��ԩ���1����G�=��W)5(��뫔X,���r98֞|2�Z�����kf��h3&i��c�5�Dc�#f��c��{̒{1m׀�k^Z�R�~�@�T5٢�/��f��+�k�c���%bVBǂ:���!(�f%�  �X�O�sN^]k5z�¾X��Ű��ŭ�m�_��U*��Jg�# <eʔ�6G�]��� Y���:f��w��,RC�p��	��e+_�׿�����7�NW^u����#�V�
Ŋƍ~��;	MjT*�$=�h<��|Ü�gBW�]'�I6>�1��6�������c��ٳA:h���0������y,���k�����Ͽ�Ug������W%pcP�����m�v� QO��X�<<v�&��M�`�<,?�-���J�.���~�(�_�\}�TNk�:w���`a    IDAT���G9�2I���ӧ' �#�����h?�7+��u
pf�%�G��q��w�z��N��A1�/�õ���0|W��Y���>�L�G.��ٙ�vN<v�����/y>���hVIs�\���y�r����FUK{hs[F�7�U(eB\=	��Y���5�xLHb�y%s=a�ۚ	�x{�qb�'� x��s�W~����&ĸ-q|�.aGG�*u��=氉'�l��|H�pt�qg��@v��$aN�p�Z�[���yW��5�2r��q�M%~o
Z˄����Ӫ���{�{���õ�����K+W�5}���jR��S�.'v9�ܙ�2irȶÑ��+MR��zW�����'C���svtt|�dlj��JaG��?�M�TiKIQ����n��ğ����{K_�)���[]��?�;�lyv5��kp�s�U�\|��������;�l���=nG�G������#�RW�f�]��[ޯ���%$cY����?��C&����N��:KeRɶ����Y��ɞn�i�1	ۙ>n��\�w��-��o�I���N�5�����keҙ�ϟ��2���5��d@�=�`K������x��44�w�"���3�p�2 �ٕ��X[��9�v����Z��Ԝ��iݚ?�sO�͟�Z��f=��Z�:�*ut7��\�t]6DI�7s��2E�
ay V@���ϔ���U]�>������|�eb�-R�L�d"ZM��[/r�N�-������F�����{0X��D�Ɇ��ҽ�1����}�xy ���緅�mӇ�a��`�����k8�$)+��|�2-Z�/��lӨ��n���{ީ*���G?����s��P�k>z��:�x��;�9�TnT]&�j%?(�������w��П�o;�I}���n���`���~o�mw_q�qSV�H�����τuk����0�R3a2� u$K$5|c;�iz���I��c�k�٫�s��wtv�Z�+N{�D�퍼l�
f��ک��\0Zw�y��9�h�^եw�~�z�-*T����<g��v�R�l0q*3�{Ad��3�-�[*��>��I�c hIo���m�3h��kGA�(�[��=F�w�~}�m �5���c���0�$S���{�!A8�pU����\m_���f�ܺ7����P18W�t�-\𠺻6ktKU���A���ܺQso����ȟ���[���iǩ��M�l&T%�M��Lp1�ZSA-�>>�d�� k?��$�^`̾��� ��cRi|�%�߻�ۮ�8a����q��Z&ӥ�M���۲WS|;�\/� ;�l��m=��' ^��p͆m��M���%��i�l,�t�N]m=����5a����懪m+W���PGw���z���^s��:[GN=J�䒌�
��w\��cOa�d�0ch���v�z:���Y�1���b��$}
��m���jp3��(ÔR���H���X�v���X�I�h�����HQ��=~{�E��ķ9H�v�r[�U���}���ѮQ�Ӻ��K5}��նi����&�ት:���u�e��ɓ�ΕU���r��j�8$��i7C���\r���;I��w�U����\�w̘Ì�EcsD6���=��s�a�6|�,�ݖc&L5@���\R��*���!�������pd�'*���+5x#(µ;#���|;WܞT�*�L����-�d˪��K�W����?Ձ�ї������?-�E�Fm�)U(:Bzr:2َ9�U��]ׅ��v�����`��̒Wt�P෽ ����''��&�W�����@̴������>��)���`~��]�Y�4i(�p,���� ��m�  �~�˖/��C]��4�Y�e�e:������������i��u�'g��#�R���i�V.���	T�2�؜8T;�s�:�#��c�F���Y&�h؄�Q�����xf0�S�{�����{�U�
�G^v�!�Z�,h��<��-a�N@8�K���[���!����aa�����l��ST&5�N� \���h�|^�öG�ap�a@!�`:�'e�舸T�A����wv���/WJ���+>r��Œ�����>���*����@u��}g���=^�<!4�`��5�9b�I�kn�[�q�$v�����@oi�P l�ؾ�a��Sj`�P�P���^����P6��Ȯ���؄��M@�H���՟\SJ)b�۽0DK�6�C�;��[����2GP[�[�\���657V4�+u�'+��~��g�������h��>v����T��Ov�	�l���0�0°�F��1�M�i͵�(f�: ��h�^��:��E0������7��7�����n�͙3��a-�~�U7�ۆ�{:�c��؄�J��l]F�[���Ïu:YU�0�Pi�0'������c����fwꩧ�z���8���/��{�e9��.�f�\��A�+�VL8SV�g��x�'�<y/u�!��˨�/k�ڂ���~�wfƣ�-�}�{���p�J=IȌm�M�!A2������w[�l���@x�I8�c���?`�j���qt�6����Ȃ��0���j�^-�m�{�/�dk��|3��(��o���n3~mӏ�@���y$�m�0����� z"��3�&�
;T,x��*���PԜ�.׌�*�+�����K��ǧ�h�����_�C4ԏR�@�U.�Sjm�1�����k�;���di�=䍲d����k��%a��l6���v�'�x��8�����${�Q�2�I?v�]s��퍦^��I�oZ�  �� �M� �����~�Lc�� �m*�6��@t��T�uvc����1w������c�=v��&�	so�f΀�%�\���U��Ù)J�M��{�Ǝ͉ݗq�Z�g�yI]x�:�R��T(R�>]o<����	�
��bZ}D��c��VL�wB�fǓ�f�m0�G0���1(hl��k~(��\�õj�G& 80VE��D�b�ۧ1���� ��18ԫv1��0��b^�z���_��ݪ�/��[.�y��b�S�,��ܢ��Ps�x
�r5��b��+µD��?�]�&��5YФ!��*8�\v҆�T�F4z��9��=�zꩾ�,��e���]
»mZ��9�y,NK�I�����3�l���z��a�"i���A�1x�#V����g��q�V/6�H���/���?�τ{�U	[ }�_[� ��N�@��1{7ͬ�w�*�jk_�Ɔ�TI
MW+9��x���o�ӓUUuJg�rw�6Y�nPkx�I�ϖW����n�֞X��)_
�℥;3)`xXM��JbL�H> �x�����g��6Ɩ��P&�>U�8��!V�X�ֲ��VD�1�}��'�%���,�Ύп��+~Nm�ĹB�կ
a�������F�]ñuu9
� �*�ej�x"��{�����I)��λ%� �O� �-�^��ܷ��\��I,ט�$~�$���t~0p��P��$���(̍�8���uu���~��}�qe�%K�����:���IS�0����j�(j���C�\����L�m�R*�jjjs��ȩ2N����\gW�g���ȁ0S�����TfK���Ȅ���P��Nv����ga'��  �`	c��M��p.�I��aA�e���q�]�L�:u�v[>��O��v̓�
��2�Q�(�?z�({�њv��Z�z�V�\h���=z�Z�^i���st�ݖ]�΃��`�l�	�bOfu��y��a~FV��7�����s�;6wl�eu���O��Z�v�Te�����ƌ�C�ֵ�R�*+5�Q=��{ϰ��{���ޤ���'O�؞h[ؾ��l)~@mY�aI:vb�J��!^�.I��e�"���8&nG�����&��+�)t�A�� �j�'wr�d`�a=\{7:L�c;�(��bU
q���`�b��$B���6�j�� Ό3#c��MS��'��"c�&�<b�N�p뢄����2�<qó`!������_�O|��8����6?,5f�-q���/*p/z�L�Ֆ
_�s��U��������=�+��6��o?�Xجa�(�D�ӄ��e���w��ή���Mx�Nz��zݞ�W&S�8��qT,�o	�����K�ro^0Q�a����wt����;� ��Ny�P"ֹ	���Ш�M ��/��!��x1��&X��6��'�%!ʢ��� ¹�G���k��'�]�`K�+0a�C���#���w���`����/���\~X `��:�4���J������}��U��a2�m��0-Pi��b���_���m��<�`Vm �-�R*t�d��*;C y]]�@����=U��/{�'gUvf�i[S6��:1�CH!�PU:�ˇ�AA �PE�E��B	5�Jo"Z�	���u�;��y�ݛ1����_���o7�3o����<�Γ\�e�!1	����Xc���J\�?���V��/�9�M�;G߳EwY)̼6�n�1�YW��ݯ�Ɯ'����8Oĉx�|l���1�
�LB��.��m
����A�o9��Ka�M-�7ӓ�GI�1aס���\���}�SW`��-"��.ס�Y]�J�	Yݫ|\��/.\ǒ�e�� $�]�u%qL�����qt��Ɉ;6@Ι����(�����g���Y�q���f�v������"�#�qEr�������ΊAXI	*r.����f���?s�!, �8�	�-�;�WX�p��o��Ƶ��Vj�7g�IsĀ�"8�����s�_~���٧���H���xI�^x��;��Q��Ր�9�9�?��!+��G�l�3*�E&f�E?��n�����OħL�p�p���[R��Ƅ���1��n�0l��x��iX0!2�\����ׁF��������:o���τe������K�������O-��|4��b��G�i�#� �͍`��)�x�|���4�2���cv��B�"K�@�A�<�aw���d�b�n��i�W(tXk���K;��%׽�Mhg��bN���9q1;���'&�	Xp�l���Ĵ���F��3y�v�r�#7Q��h����u�����x~�)����-��Il��t���p��Y�]���������M\~^��B!�O���g��j^��KznceׇRU<�����a5:�qH<����:	ܦ"�s�p�A`/vk��W��6k1o��;�2�x%A�[�S	�k������\_�by#����o!,��@R�Ϛ���	ekκ/��B�4��phqR��&K=�s��:�����&��_��5�y�d�Č]w�Ç7}VSY	���6,�B5���O�In�$���)S���^��)(�㱻ϟ8�Ǜm���e����[q���o�gќ[	�4��p5���H���^y�v5..�^����T�����e��鲛�c�=��6����(�����o��Ád9�	d�t�qqˣ�����R焍!��k����s�Q���B.��H��#W4d���>Y<G`󻓁v��0���um��i�S�Dt���a�d��N�E&78����Kf#UE�t��X
�{oQw00N)96L6K0��"�O�}3V�\�@�G)��~o9�c��e����<��F������T�0�D��ɘe��N������ۏ6�U�Ϧ❖Y��j�MQ�3�Pf���-�)�h�ùm�<�4U޳���˷��E��7�>�6T�"!�yw�&��O@��κ�g�I�):s��Yleˍ�)���E�`�M±�~�3am���ֱ���e	
�����,(ֆ\˳|�`�e��6Dm-�J�_Ѱ�b�b�$f�6LwL�i��~�3�u�Lc$�<���������_}�J�e�,�����7�4���0ٽF��׿�9�;��8��2�}Sfu��0��X�΋.��na����?����	��m[(9�{�9�s����"2!	�LI��JiBp7�JoaýѣG[�w�)�y�lxI� 566b�ԩ֝�裏ƨQ�p�W�.��ó��egJ�)?X���t��{�>�+�Φm�p��Yh��G��6cCe�![��P^�![be�N�pq�j Д�C��T�0�����C)ӈ�P(f�;{����,Í�kC $��������9b^�!$�Vf<��-����6c<C.H���]��.����\�%Ky��(����N��� eN��D�{<F�Dc�H;�sa���%���P@2�p�8S�MvW���L�������ܡQ4gn�����댚�Mn��p�?O&�+�ȟ��ʲ�9�'.ŀ�Y^?磫0��g�(_3�Y�,��ٹ2�Kõ�2�J�S�'����2i�*Y�Ry8IT"�d�o��ZfcXB,pL���'l}�Q��䇡��m��E,p#d����#95c�2�aS���8����ǒ���޸֙��O���� �,�ʉWd�>� ���_1bw\x��?�V�d�Esn#s�qm3|+|���������3?C�fe�Ձ�d�2�������"���3L�rPi^h�A�t�;�hM29�P���n�B���k�ΐF(���@g>v�<� \D<Z�[��B&�;�4f$@L��bY�$�vg���AT�[��}����t�71�yPd%0ǂ�1�x<06l�/:�� ��W�dO%�l�fs�NB1���f+e\�u;�N�عr�	XB.OO�[5�B�͓��e8qL�\+E˱�%45-� ��<i��5�g���NOfb�����j	dy�sx9&�{w&���
��W�{�F�nFZ�Ӳy�/c�9nv�n��5\:N��-��*��(9& Vŭ�T���?�.L�t:�{~����@'5e��x����:	�1B��M~_,��9G&����|5�<��:�1:ta��� �5(;�wY}���y}��f��,T"�CaB� S����'߷�%����*������q�Ɋ	��gZ��{y=�2���;v�������UЋ��t�I.�L!ي��嗝�X,�h�x��d���z�ͭ��X�.8��n�MN8s��f�V�n��9�6#�a����}�*(��wN�{��9�xѼ!���mg�曩|�4/��n��L -b~�i-�4��N8�{Ԇɐ�ߘ����tP�RϪe������3���O���մߢ9K�vʠ]r�h"�tXz�	:�r}�R������ �@eig�9&�r#��z�������O=b�$R�u�IUaIK��/�ʹl���mns s��4��A%9�ts��qV��%��>������ NĀ>=�@o��M�,Xf�6O+�w�f4�B��%�h��ȤsH�T[��6��Ǥ�Ǆ����K`�����-���X���bsk�ѷ_O��vC�݆C�*E�cP�ˆ�����ظ�D-r�<�j�1|Ӎ�e;�ܷ6�"�!�Gj0o^#>��3����������ݕv<òsѴ�(����·hk�!��6��Z{�(�l�"R��p��7��#H��fb�%��Pz0�76�p]�76�q���Yb�N�)��%����ȜĜیJ�x��У.�|��E��QJE�:�Ut��;g!>����q��O?9���4�ݳ\:��X+��ǐ);;��<�2ea�h<���� 5t�1D����&�u#�Aa�}Y̼:�H����B͗�9s(����H�د�l�N=��M]n��E����N��K~����9�x����;����"
� 2��s�>�[3�X;��ܹ���۷�>�n�b�Q;bܸ]��?^���s�	r�#�!P0v�7����Hy����,й���h��sg�Ճ�Nu�q���������>��c���ꪫ�5�嬑�T9�:��	Z4��	�?*8��꾻�d���i�jg�0S,�A"�g� g��x�5�$c�C47��F��d�+�УgZZr�b����_`��2�L ��{���N�.z��Ҵ��uJ�(|%�d�s5ҙ���V���_,���ev�5�<�$\�\1m��	^������e�����p%��    IDAT���"_�p���}p�٧b�&k"�ʡ� �L��Eʱ�b;jkz�����^�ioʹ��h<�w ;t�egS4�B���w��Ƣ���-x���n��6���@�^Q��D�Һ؜dEz�I��)�t�U���o{��L�Q��Uᢋ�ða�!�����i��"��"JQ�o'0{V+~��3��L]��^=�8��ð��۠��N>��_o�����Ǒ�U�W߄�S���O�9zc�q�ѧ���:���ɍ,�i��X���p�ݏ��߄L��G5���ß��}z�O�!�.搨�E&]v�E��T���᷿�f�Z���1c�G������kY��B9ϹYlPfr�	���^\���ٯM�M:�	´�����YSr�If�8��~{�,Ʉ�|�}�w:�h�I<���>��S�a�� Y����$#vQ�B"�|�9����v�'|����]4kR��y[�4�6�h8=����VA� �L՘i,t��yʓ*p$�e���	~���,(A�7��gJ�
���79�ػ馛:�׃�j~�Xa�:\���,Y��c��V%GÜ�T��gc��F��i�(z�^��۸&�b���j�z�q~�r*f�`A}���8��q⏾�d"�0��L	DB:G��������<Co�5��q�Uȴ-���7�o.;U�EDb$�=Ē`B�:��96���}�M�?�*,\�A�cР^��տ�F@UMK��B���%KZ,?�mB}�����y8�?�g� dM�h�?�;�\#�|����ȤCT��@1�As[�9G�~q�p��Amu�\6�r\���У��E��I�si�riԲWU)@6E����wN�E���b�^�S�������2��t���׺���6Ī��a��-8���֜4pC���y;b,��<��zd3�9]]M��B���5ho���s���}ɮ�6ဃ��ŗ�eV_U5=��҄H����$r�fD#Z�C���_q��? �gDK	��xn��r4� 
�PU� �#yh!�E�Q|2}~���a�Bnp���5�G��/\גDW ����1˰N�3�W�R�+�>�� y�G��Z%0r��QG6K�!A�~+̑�F�ʸ~�Ƈ~ءo���������=�S��;�c�Qq�a��*�-V]*���x|�ĉҭr�	�i�?�:�2B�䌎���:s��?�~�4a: x1��#;�7$�P�T�p8J���@�T��M�j���hq't!1α��\Dw8e�H?s������y1a1hm"b�_�u�)�����z�U#�m�5� ��C*�ܹ�0����޻�n=�[�a�u��̚��u���q�DZZf���cL��.�0�����O����ת�&Ç U�B6��g]�{��+°10z�!��Wg�GC�X���2M��1x���zۍЧo�m%<�ī8�UXҔC6���5{�ګ'bذ5-�z�&L�`f�^�D�
#Gm���kP,�ha��#|:�yV�����ӱ�ޛ��g�t�^|�~2˼�[l5n<��J/'�����Ȁ�m�&���r�� �x}0�0mm-Xc���醨�AP���;����X���q���a�-7B2Z�3fᓏga����Mb�m6Š����=�Y_���C��9!�R=�f��3�����BUUm�Ux���1�3����o���,"h�9g_��S���,��"|{�m���~�T��%L�����4�J	����t�:����}n�4��t��Ym�h����5�ć=���\�Ӧ���K��l3bK����|	�ޞ�SN9��f�h�p=$P��A��Hi�_g������qq�+.~%I�좋.2y��k�5ف�ε��q��g[� �F�>]I���d/2W9��Lc&�Z��������˟~b}�+�P�Z.�b�;'N�����?cH��_L�ɶo�L���܆�=�b�}��A��5.V��r�)���r @48�*��;$w$F;P��K��?C�7��.���p��Q�9?TG;��&�AO'�"�4�d�c1��d$��`.ǃ@8Z
Odp͟.�v#6A.�Ƶ�\�{�z�L�d�l�)�8�x^k >�t6�9�44-�6}-6���N��(~�Y��������-ns�o5��c��^���b�s~~��o�ek�JF��f�����ƚ���������Ghoˡ�z���18���Чa �|�e��G5hM�bР:\s��>|]�����<���hivyc����~�t:�c�>�L_�b���
??�T|��/���)�������K����V������{����������)�DX�>������Ä��_y#^}�V�y͵{c��vŉ'� I�r��8�j�Zcu=�����м�	����x�����j����Gs ��>��Gu*�|�A2Q�T<�?;2֢C�L~7�x7/\dRĺ�Ʃ���ѣ�`�b����	���=���~솸�Hā�>�<~w�x��/�0x@_��q�w�������I��o�F{:@�*�~��4�2�ѯ�f.���G<�̋h��|���Gu �Yo}����ޯ�����t�0�v��#1�n`	K^U/�}#q�V��KVvmq�Rz�߇�0�F��ɻ����DKZ�*�Đ!j<%	&������E-�Y�_�!�.C����'̰XFr1Ȁ�r�H�D���O�֌9���1��ɶ���,̇�S��2�v�c����{���a]���29� xC���!�exژ1c�ǝ�;o������3��Fq��%�s�YҒ�뮻����4Ox<�QҲ+͉;�9��K�Y��zEX�M����&g�:�z�1��`ܸ���k���������j�`޼�h�_��O9�}0�,n����%qsƤ��8��#�����s֯���o�&5������������~���/���Q��ZD#E��.~q�9�7�?.��j\����,�b��=
�����1��٧_'��$�-d���^����0|�zx������}�a1�"Wh�O�8�]c/?������tR�)E��s~�������<s�8ӢX�aqS|o~y�D��q�����?c�� V�&��[�E���e�^�{�~
�4��#�������?���C6ğ�<��ş�̉T]\�s0f�V����qٯ�-K���ޞF���<O��T~���p�yԉX8?�T�^�6�}�I8��=1�Ïq�����g��"��2��k��췿A�Ǚ?�S�>n�z��{l�_]:��/�◗�_0�)�$��x�6��.9l8�L�Ɵ�G�"5���֐�x��̂����p��+P�Ҫ`�q5=����}�݌����s0oN����lQ ԃɄ�E L��ײOθ�y��5��Ck��K/�O<a��.�đb
�$��R�rY����$1��u��� _r�wՖ �&>������z�vN�XG"�0��5q��S��7���k��7������t�Tס�.�_���k�=��:k�i���O]3���y�^Pi�t:q"����d�,ʜ ��3��w5������w_LFN0YCF�������{Ȝ<���X�I�U؂6�Jv&O�d���:�Pl��ڶ�����>���o��C�����h�^W^�'��һ����p�i��\��	S�~�s���`�� ل���;`7�g�~��r/Z��[�������x*�)S��鍨��l�� �G�� �=�������	�͘c�o��:��ʘ��t<����=�V,�U�؊ۭ�]v��By����x��O��=�z���N�ƛ����x�Ǒ�31$Rq̟7]��{wD�$}�9�v�ݦ�&SQ��iss�V���;�'����/2�Y�Яvt�>Xc�@���?pß���y�{��:}q�O�ƀ�x����g_B6�7Y��nɒ�a�15f4��<~y�o���_���Jओ����73g�#�����
�B(�h�B}�*���H$���C��ǟ2���6�}���/r�y�������OQW�a��l��y��X���6�c��������@x���8�'G0���0��� R� �@u7�F��ƌ���M�﫮�'�q9s�1���%��rK��rDe�D��EI %�u
�ZS$I���A�c+�%�����Ep$8��O��"�����~%FWP�,*��H��K�@[�K���~֡!�f�C�|�U$)�b��.���w;�?���\�H:�k�^���*K[�e��H�e0{�\�1�/e�H㵐�04�L���ed����l:?�L�p��Z���~�;�ŸH���5N3�������mI!+zМ.��K,D2JW�+&,JfN' �0Lۍ���ią�[ٌ��̌�\��<둘�a���;�Xlfu*�	'����ej.j-�!��X*ЊR��
�B�5ep�ͷڦ�H�=��[l����e�!��^��
%;�'�mv����cūo��X#Fl�q;�E]}5r�64�����X�Z8Ya�#H0�-���>�*��y�;dm~�Av_�7$��%�d,i�0�!�K�����0��|�-6Gz���~��dN��C1����JAU��Rֱ�\S�����c���a�=v��^
]]�\9�9�k�g��h�T5�z�I<��S(3Xw�5q���G]��7�7��_�A��L������,bL����%QW_�}���bNU�&)�N��u��IV�"��a��&���x���P]�n{C�1p��I�NQ�Gl���N�P�#_hCMm�eT>�̳x�o/x�i��ɣ���י�]}Wk_����(aE������H�3}G5UH���nSK4��G �c�ǣ��r��7�҄�Yeg2i��(7^j�����r�A)�H�}�9���[C�Ȅ�͙�F���ie3y$Kq˲bg��F��vێ�@tj'�%\��+Y�?�+Qb:!���ܝ�\`.vҥi���;��LX���|i���o?|�;߱z�<�@W�&���,'�o��{����|&�0M�]v�	#G���{�P���
�X���1�ic��.7�x�̥���ȣG�:��T;0M���Q���j-0v3Ӟş�x5�45�Yz�!�c�M6�D�D��ô�(�j{{K$��G�0�H�}�Nśo�D��a����hooEmM�|ȸk�YSRr������g�J��Ͼ���z޲��[-x-�r�������L�̤a�X�u�]k}�^=�C�ydŁ�ģU���N�!��1��af.d�����m�[>z�Hs~Qv1'pZ1�L���X2�x�������G�X$e���\3jj"V2'u�z��Z�03���]�[n�dCF�q�!Xk��(�]-�|ԅp�r!Xl(ɢ6��A[&�|���w��=��M7�L���8b�h�)茲�����H%��w�Y�)NX��-����kM-;��s���Zת)�26]���|�2�8~�R�E�$W�B�N}�׵�n%g���H�k��GC����s���;�k�3,�8Gi��^��p2����/>�[���c��Q*o��jy�ąQۍ��oiT��7u]� oȘF�d���E�I��aLa&x���f�>c��-�,���O3qȄ��T����yv�[�ʿWFX���06��λ����0[��w3�ъM�ooO{��2��wϾ8�cгW5r��9IYt�]��ɞdɽ�T��I����Cs���r46�d�����43��h9���&�4���g�ex����B�؆v�	;�ݫ��ێR��[X�n��W���W_�#�<jbk���q�Mb�vc�>�V�%��/:��y�����OV�&!%*��&A��2� ��;�[/&��z��������0v�]Q
�`� 7�(#,��Ӳ�-6�.���yx
�b묵6�8�H�V��4�H�<��}۞�Uch��'0g�b�1�n�e0D�����A�LCfZo�Y�ш���x�Ld`z4"hko�=�M����7��cϽ��[wT^3�>t���8w�RLRJ �i���?�g�}��	slx��#{f_�W���E�$�I�fh]�؈Պ\�s[�1���,�L�Y�$�>�E��A-�?q��@,�:��tApϹ���ne�C�?k�~?�T�ό^[�b,���ײ�gRv��0U<F ��M3Ώ�I�X�U;b%S��)b�0�$�i���IK�`� ���d�(myUO�/s|MM&��Qc��.��B����VኺS�'x�nU>x��0�d����w,�{�P�f��M��S�*���b,�l:���x5��̷B���{6�h0ق)��x3��ƺ\�6,PJ���x�W�۱�.���ݝ? ��5W��^JaWq�����w���GQ,�0x�z��P]Ͱ%��:pP��Jt^:	f�������Q��Q�C=ܬ)�"��X�,�+�t�v�w�]6�8�;�;v�
�@b��<�Fj��]�&^<��sx���a���z8p�Cѳ��B��`	",�hŜ�BM����1k�BL���z$r�Vt��/�"P���]��8u�b`R����<tޚ�������`�-G�gى,q�R�yj��t�C5)�z�	<�<#���)��V7��>h+���X�"C|8J�
  VY�hԞ�"0��S�	��Ĭ}�/�*�Q%r.�2�a�_B�y��R3!3�M2z��/��Ej��E���w1dW�fk����!���x�*�n��\Ԅ�g�6���;Ժr| �������k2'@ǈ#��.;u�׸�0k����\55�V;���>�t&�k�ջh����j���!�Rk��z�e�o�|7�)��X��s�!��Łi�g����E�$&e��5&����:�_�p \(�1v���N�:�-���5�\Y���_���NE.ߊ!��G�J]�BV�rV�c���X91~������N�Z� ��p��n�~J�r��e��E1���]�h)��v�;�0�
Њ0RD�M�D ,3EV���A{�ox��Q���zb�}@C��(�Pv ��v��Jr,�4{�|�1�.4��X����׊�S��2�T�t�rW���@ A�<x7�}w�""�b��lC+�K]�9S���u�ؼe�&"x����⋯�>z�,%s�r��^��u�g-'<׺�[��t�D�H)���"�:�i�������*0}]����~W�2Y�d¿��/~ԭrİ��f��ٓ��i2�@�@���m��紜�dҨ����	\��:�/O���f#���Xd{d����T�e�����oO8�L�%���"";ﴃ��O�r�٬�?�0�'�|��������'N:�x$R���E2�@&�C"Ve��`,w���D�=�o��g�GU���{ ��a)�"� �O�"�Z��=�-�*�?��|�D�El��6�c�q��zư�Te0�����xO<�(ҙfl��z����0�.�qԚ�������Ł�o�h֝���_�>���՚����u�ݹr�1L�4	���9'�����a���23�1�HH	B ��� %��ګx�ѧ,Ds���Ł��L� �M���+0�w�:{�,�:�6��6��G=�w?c`ٴ�$�"f�k5����x�-���{��p��6nl���	+��Jo&aD	�L�ȣTt�V9FO}��K&���bC���~��0֊�$U"\>;����h����ҤŬ�m����9߉1���o�r�y��K.���
~�g�{-�q�@�J�\� a %k�����H%hT�?`�@�Kf��KS������J��C�J�_��<Mؿ7j�����:��KC
������P��*�;�}�|���"��{��O�z,2�8k�DV�>�:چ%.>�����rf�j4)�a~Æu:)��Z�h	�@I�d�-�G{o���Uy1jv�aL�ȶ��:�߲�G]8���7^�3�<��v��z���}͂".]�[k�d�%���0=�}Ѣ���Y���F�:�k1E��[LK3"��P.IF]\��    IDATO�ܴi�%���{�յ(���61i���0.�*av���x���:���?�PTW�L
	�1�y�e.l"����3q뤛��i�1��?C�Ym-��y��PaW��Pb='�����R[U2eN�-�����:qƨc�ni���qh9�C�ԩ���^� a����X��^_���V������'>P�v�S$7?��O��O:�W8��|g�_U��Ap�������[�"+�Za��3&��c�Ǆ�@�L;�����r}g��8�J�
�����:��v$�I+9��c���ϛL���X;c�]�2	���+��և�&�5It����~�L��\CC_k�Ds�Be�.vR���R�|��b�	sF�>�N|1s�1�C:n���0z�XP���ddtƱ6��g����cx���p�[c�]wq H3Z=�:c��;�i�/��"�y�)��6a�����|wo����i�ńs�E	�w:��;&̤��o���fs��0x�Z��v́��`�\j�cA����`�;����v��Q��F�n�:�:4����x�W_S~�tu�Ї|� �ץ�%#N����Ps�����?~��{�/h�Ƞ���m���R��G�U�c�>Kf��1&v�=���!��[��-�ڼ����\��I,��4~
"�pK�>�����_�waiƄ��L�(�b�7 ���^O�����F��'�`�����U�
��b�>�乕����?��n�ދg2Dm c@��� l�˝'*w
޴
t�������BVV�~
�gU�A������u�T���d��׹x"Țcs��#)����@`�<g��aޙ��y띗��o�vۍDM�7�"�;��,یBgqmV$���v����|��6����0�5��$���='im�K$�� |{�[���f���κ�p����$A&�Yh�����:l�����&��ʭe�/F-8J� ��:�!�����|�m�PS�[l6���6p)WsN��~o;Ν�ޙf��'�����:��b���(Wi��R���@&��O>6g(+�54�[lf�4	�iv��|�"�ո���z���4�୷�FS���l�a�ӷ�1ב$�u]Fl�c�W��ioǻ��f��߃�\Á|YEp]��Ȯ�5#n����������ˌ�܃0�,"ʝ}	����}��+�o��6�Ë"�b�>�7������w���>+�\j��	&�ԭ �ى?ԫq��u��1%{���s-�����v���)Mƿ�=Q�j}^Y2~ڡ��ΤA��͔�8�?9:ƃ1�1.�"�S���5��+6�����bE}���L�B�ь�l�����v��&:�Lg�p(&-�>`�VTUV>,A�=SDUu�����QưMҊ)����k[ښ]�*5���3M\' 깱:�cîȓ
�3^����<��	�S�����0��=,�M)�oG,H!
6��Xl����խ���uD��@�E6�⅝%��*�=�v�p��+shl��64�%Y�k�i�a�."t�#y�-WQ~?�X��Y��=;�7Yk4��k�8vڣ����
�	�s9�9�)WX)� mmtF�.��"C�z���;V���Qu��#X�Y������8��J�}�O�ӷ�eY����O������ar6g+��D��Uµ�V
Fu�7����\{#G�+���+e���H��i��X��~�Y	��_���vl�C
�r^}�cuG����r�t�q�c��/��u�y��Gz���g:�4K;j��v�0����`�|�g�H	7�.j�	�e'�R���s���˭(���R��Ҟ;�
�w� P�K�"��pz�����d�K�#W��%���ʛC��7�-US�w1͝��ܚ�l�c[���p|e�	��u-]�}W1��h����z�����]!a
Q(r�3�2��QZ��}�\y߹���y�h4���	N�V&LM��a�X�av��!@��I#S]z�;k,}}�����^Y dE���Ү��U�B,��n�:�@��emB�{>�𿿬��i���X6w�������0�<�\|J���;�ry�]�.!�+3_*�ϲ�>�,Ӻ������蚻����o�g��i��@�oS}~��|�h���g�>��j|�N��RZ���τ�ͼ���:zy L�/\� �O>1_]���R�v�m���[�B�&O,�ں���\+�,|���	��]�ݲ��r2��}���X�;�騩�'��D�s��%�2��د��WW����_����9���|�>�?s��k<T���-P�wĈ�ch��y%�O�c���W�|�&|�y�حs��3o���6���4�r�����)��O o� ���=|�lK��nQ-�~�&�׽��YWLjy��
<W����8�;�oو�빗'��^�2?�u���l(��X�s�Y[%t5?���|C�,�T9����D�#T�M�$�h�?ʟG�/!�X�Y�ڴ?g���R��{�'u+3m��B�	��Z�</��k+5-$1�J�݊��R��`�;�����}C���et$��e��������|Y������q}r�U�Sy���돕�/�[lV?�?��_��+��O�8珈���	l�3�������
9��F��KN��R�,��s��I��֑�a�i%�w�7������.e�q��ޮ�F��Q�
C|����Vf��_���W�����W͕��(��sU]���"��b~0�@T���7���z��������r���խ��g�v�X��q��ܭ=�6��C�/�u{}�u��@�2�XN�P0�d`0�LqxLd��L�L�����Ϝ+M3��W5�W�����Y޽�*��e�mE��U�~oY�te����o�g�.��{�:��M�n�cޏb��STWm��L�+�%�7Wa�:)�H�2���,@ƚ�Y#|Sނ/i�|�b�H&|�E��[Ax��g�װ�Iu��m±�Ӏ���5�ʾ1/~��@i��a�(�]�|��T9〱�o�5e9pl����dG���T0^ނ�	�������u�/ouu��:��]]��t�	��*k��ݿ�wI�Xs�䎅���&��}֩a3O&�̤�^ͻxh?�B�	��|d!%f/�>_�G&P3��UӘ2�^s<��=զ�@x�E]��n�MN8s���f�R�k�jQq��V ��1�����f�a���V{�`�!��y&o�i��Q����,+Ț�
#Q;i�]u��]�۳Xw%V�g7��.��O�0������*�no�����#�F@&?;�����	�lgĵOF��cc�I��8C�&�BE�+,�E�`�`�5��B���bb�AbI<#N�K<�=U�����y ~�\�-�ܲ��<�֎��S7�;o�M=�V�PB*�B1��v�l�]w�Śpr� �U�y�BJxAܱH�Y��Ay��g��B��~rg#��L�gђ�>��w��3����*w)$�������J㑘��v�4��`����X=�� ��{��h�����@J�5u�T�u�YV�N���׋��'���'�"�Na{5Ue�3�?y�-{b� �?Or�k�q��*D��)&L�^v�i�4̟w#��D��
1�1z��ǖ�l�-�9VJY�m?|�]�D.��7�Ϋ�9�2�Ѹ�H�э�{�<�䯹�c���ؓ��m���G�?��J�p�k�M�_;uV�m�����-��.��<�1b�=����=(Y���+�4FK"'�� I�H�j����*J����ĺ�C��J��CI���5�᷑H$O>���O�V&��N:�i������0g=��F��9���z�V�a�м�	o����=�
��0�P?��7�B*d���s��hj3ou����47�ݔ�̎�,���&8���oM���P������zV���~H�Ȅ�;�<�)S���W^1��l�w4)����aGr��[}�X�/�j��v����e�[�8�7��|Q$�$�dƊ.� �A�}���� �gќ��m��Yky�]����i�ѧ���[vA*7I�+�W��5��;1ی����R5xj��A:��#�	Ҫ%L遍?�P�;�\~�pw�����3���#��� ʾ��%�p���Q�$��_�����2�
/��0t�P+JФ�K�!�v�������}=e�w(cЂg�]2r�����ly����� ܻq��#�m�b��Sb������Ǉ��?��#��7�~����y�d�܁�w�d���Ȇ))(�[�+�Ѥ'��l�i��&[%qP���Saq|�����X=��#�g���;�Зv�n�ă���o�%���('���M�GL혟q�Y�
;#vH��(W(m��S^��x6y�d�)|
�0���<��s���[/�2��Bǜi�o�/�o�Z��B	}k�X�چ<�ק�7w+^$���YQyi,�$��N�⋀��3�4�=��y;��q �w+��������d�qJ�)��|��� w���ek�gW����׎ q�k}�]v1ٓ��H���I��7#���0?O�ψ�A��Ad�����^)��O,cH-ϧ�3C�Ȉ� ��N�9A8�M�����#F,�2��%�il�!Ѷh/���N����/��q��oܕ(^��r�� i��	e��)�[�k#G�4`e0��;��q�g1}o<�!��t�I־��=w8�<�����`��Ϫߙ��Y6rU�q�qW���pHA=�@K�E�� ��{v��������"��ȓ-��s��̗���@�Cď�%&n����o�u���������ގ���b�L��s�9��
��ƃ�̽!ֲp;�`���c�=�������g��5O���]���y3r�|. �勃�}�-l� {�-����;������8h4'�B����կ~�O?��cpy����ᦩ�����.���R��Z�l�cA��ˮ30�Ė���x�ڳ�;5�/6h\�� �M���u�*��+CBW6qey��5O���^{YtgX+Ca�W���β�ӧ���B�����a�S��B+�@���
'�J��$~�	�%q��=d��AxqӒr��A4r���N�V9�q���ϻ�>�ގ!jl�2b�m��|���2>���fk����x#�q��͟8��f���r���;:2�)����8�ṣ��[����}_q��q����zt���0�l��;&��^w�H�QvSP1qW�[�r�B��Y/�Q �=%��`�)�篁/7�2�_��LE��s]o��&8ꨣ��&����QF�����]E��u�]�鐣����'Ű5ʜ���v��9AX	�Hi}�w&�͙7���,����Ϛx�O�n9���5�1קq&�5F�!��n��6�g���ן3&LM�J\�㖄A@U��&�@���]L@��ɠiV�'��� ��F�X`f�q0��@�m~���|2a�t�	�Ond�����pvt�X��B�t�DZ����Q	�r6̐����	��-���?wk�OY���������Ĉu�w�u@�r���&h0B���O�x�	�%��\�#\�N^-iʝq%�������!���Cak������9G����.�J�XL�x�ğvktkG�Y<떪�f���^d���18`L��m|:�S�J�1a^w��yy��&rGVlވ#�D�A����$�g��[o�մ���ƍC�^����<�b�<��/1�Ck3S.��q�h�%O��w��d�aW{�͌��	I���6���������_�{)�m97�^^%D}�+�j�U��/���c�=f�!��W�ċ�������R�$�aZ��I	hI iE�	����+�1;�x%�q��M�L���#A>�����v���3�l�s[�y�H��Hk��#�8����7_7&LV��߿Gș�U��w��F
B	��9m�4�9�q?��Qf޸^*�̸=?/��/��$`70}�~�{�i�1���v�i��[	�l]����>i�)�ɰ��Z����uG�g���(�9��Z]�]׷,�^�����ծ���8��LΤ5L��+��{�a�7-d:��������ә���/j�T�A�O�ϑ�1�B �02kFy1e�5��q-D���	�׽!j������ϟs{u{�1a֎�]��~�j����!Ӟ5�w,�0���
j�@J���\m$�=�`�.F���Xڎ��aFI��/A��#$�|P4T�G�+��Z2�=�uK��O������d3���b۩W�2;���_�u��d�����XU#  ����-"K˻>��I ��</�</#�ԉG;��~(�Y��zU�	�0�	Ԏ������<.�%��\"p$yLS�̡R��5�>f��~��b����h$:y���u+fg�>?�T�K�
#a� ��$��;`�m7Ō/>�������f7B�T��2R��<�
��	�a��<yS�y��J���Ȧ�"?�~�̕��#��PcE��j�	���;`e�x���.�l9��٥^�Ć	��Bgw[�-Hf;�կ�#�*G@ �*������Yl�Iv�'d�
����U��N�{�)��}衇h�5~v�t\�W>(���+�e��~��_��&��A\2"���0U�̚�wx<5%�����ǟڭ �s��̺���UB1(��1d�:�k�=PSW������wA`���0��@%�̙!&|��ݎ@;v�X{���u��-z��yY;����2�H�2 ��բ��Z�.�
��9C��|��~�����׊��� ������,���_u~����X�3���yN����ԕ5�c+ոJY��{t�}��Cɒk��	����,"�u^�{&`�ES��ڣ�I����}���x#���)�-w9���\�`�*�^������U�x,�(�B��[�w�}�8o�O��n��!�F�q x�����(Cpp1AmE�9��E��jIȾ��:Қy��c����K.����_<_��@��&P��(˲��(r�J����VԤ�(�ӈ���C	���x4�I��A��kH�CD�Id���X�C�E#�J:3&�/Z�q%��Ǘ�Rc���{��eW^����9D��k���/���l�%���&&?�0C5S��<�N^�B�����ɱ�qP'��b9u�<����9�8Q-:9p�hx,��j���gxG��+IH�m�13gy�^����]�@�/E�_�-eUE"-���|1`ݏ����4oI~�,�"Q�X{�n�߅ߣ��`��c^����sI����4?Ck����� ����Ngc��M�_� N)��=�e	0���%��!G�|S�6�(,Z����<_�a4�<aw;f���|fT�����r�G.�E�=��C1f���drvQ�UGXT "vJ�7Á�.� k�&����R����m�8��=�<���ѣ�L�����"�'k�æ�,(;�J�!�L �s΋du�]{-$�r�6��@��A�G��C,��T, f�='i�a�)`$�L�5(�R#	�"q���b��/���D��q:�GhN;&�tj�9?R�c(p)?���
,����n1��k% ��Zl��$�Ȝ��;H��.�w8�A_תI,�����ܼ_��.��k��<�ǿk����Y�k3X����k�����>��L�x�zx\���������� �����5�s���9�
�d4��|�o���ᤵ�Gh�&'`�>�(mꚣ���_�y:�&L�`>'1k��X��n˪#(��h��}2
�X���#��$�3=�_�Q�xn���11L��1�U�Ԅ�Q�gFK�H�!��fQ��QU�¨�Fc�-���4�$-B�!x��#L &�gf�2�v7�؊���:������.�IC�&�r����	;.�'�MdO����ۻ���^�߷J�,b����kò    IDATA1ӌ�TD,( d+ˠ+ҝ�n4@�!ϱ���g�%̚=O=���'J�gsK'y��X�A���;ݓ��d>;Hs��4bv>��ܠ��yl?Xݟ�Z�:������E�+pҵ�!�ϼ䑖�������siQ�㦅�MC��B �3>ȋ��z�U��[<��z)�Ō���i�����|K���;����9 ������_�;Z�*1@B��?��dA�ei�iMi���~�ZW=?րa8�ψ��+c��\</}G��~�9�YqQo�~�$LY���y�_���)�L���\�VF]�4ymd��+�?��12��f mR�#�s	�t+6�܂�'�ȧG!Z�DJQD����@8Dd�Æmj^Fޤ���<��� ��:�-(�s�%V8�v]NID&e���������gQO��gpZ�2y,d�l/�#UUg�m���5����>j�QD�,b�,g}�|�bD�A�|�-GȀɎ��A1���$�u��{к�*J1̞3�b�h��	�st��\�߹�k���$WcC�6mP81C�r��g��r��4�Z�3��bx��Km��p�	$C��\2�x�ƼV�u���d���g��|����Q�h:�3c]��bi���,&6-0��ߠ���%	F�6�y]<�����1jc�t��_�9I����6$_,_l�1�$22�Y�׿�u�s����Z/��R3�5F���/�[QQ�L�o�]�$���J\�u1����\���c�g���f˵ 4��q�2(1�:9	²��L9&�I��aj�G���ɖA�-�)Gt?�_���5����H��cH����e��0o�L��7����M0	�d�d�
�֮�3�b�.ԎD;���Ŕ�(��w��9��N��"�Cј�-���nM*���$�!baI�?A�u!�p�B>�agA���l4�d}��]��a�D�%��ېˤQW宭-�-gй<<�G���z������)U\��@W�T~���h�*�G�\�W�'�z�o ǌ��.m¾i��A�����'  �3bt�~��Ѧ�"ޛ������R���6+͛J�Gs��)�S�S����޵�h��f�w	��}�XkbYSX?#�Q&�/���;ǘ����܌8b̫��y�U�r�9
@}k��'�+
��:#���ճ��7�a��w�'��K����l��*�Z��z�x�}�!�����ƨʣ�<���K��DC��嚟�&�{Ձ��ųn�J7���g=�"3�J(9�9k�IMX )-�T^��L�@@9�r����Ap�5(��q��C���~�>''���ٺ�I�'"�DY�ǙjټC2ՓN8���,�����y�GrHF��GX�����&E�"U���G��C�A� ���g�m�H.��]{%��i)p�8�b��G1+���.����)9F�?�	j��y�1�D@����5���O�_ % �=��@Z�����{�b��"y�b�bx�C� 4|KJ��a���MJL�x�t�bX:���Jc�U:�ym�E)psSVKG(�')H�բ׳�����32�}��e��� L f��ƘL�a��/��Ȣb� �0?�Dd�g��dº����>����R!�3�j���H����Ot����";ڀ�1K=W�O@��#1�H$r�����n�#�ַq��5��ѥHj�t��sH��h-��J(�d:�db)(wPj��G@�7?5Ȋ��3M��	[��	�<f< _�^:��qmU
'��X���!(��D��>F���R�H�@8w����W�"����*����ǀ����&j0{N����6c�,���uf�UN����1����K���D��4`91�zeJ�C�����O�e-Mx��򀋭qb��3�$h�Y�(�c�͚�D��1�{qI���6�JYC�$�3�g�'SK����(V� �����3�ߡ�Y�RR�\��`l��DF�y/=R�K�b��d����\��~�z˓���x�rF�=锲$%}h}�F7?K}���63�a(�֒,��7�	��#AX�Cf}#2e�u@X���!ه��¼VE�p�@+�����z��X5�-��{�UVI�M��'vo�9�	�
s�)=���9�	�YR[��<a������;b�S�����0�]�L����vP���|M�Mz��vYǜ]�xf���֣�͵����5�Oŀ|R���E�0�m��wA��;s:��F�(
�8r�v �}dP$k���9���;��ڌ�:gfs4��"�ܽ���J(Q�F�C�z��ۏ�������q�@I��u�x�g3>�3}K7�Gm
��٬ed��0rYT���1����v0�e1b�9��tJ���'k����u7���6b���X4[� ���,�5p1hް+�*IKڈb�� t����dN�\�!��y)j@�7��	�f.V�{�Kf�Sg	�Z�҅+Mf�:5S��� ���6TW��*�z��n$6��9�Pda�Mv&���̈� O<��������W����xɊd�e"�2���j`�0&k��W]uUG%2����,��{d��X����ؖ,bޓ�
��0a~VdClT2�oai�hu�)ʗ/���z�Y�֗|�o>i�����]���~���lp�E3o�˷�	3�@XrS����v�x����Â�l3q�0���C]*@�Ў�X4�S�ZQQhkrR�̲� -�56����꾨oX�d҅ �-�-�݄L��h2���3�dA,�W۸HG_A���=)sđ�߷�*W_m)�A����j������'�����Ҏ���(����!�T}�r�T���͆�[v��MNV�z!� N�H��1c�
{~I�P1�
�z�.�b���A'3W��En<b6��8�`Դ�V���E2�� ɾ�D-�gs��|-�s��&��Z�~��YM�m,0Es��O�\9En�ǝD�����;��$�Bi���"�K a>�L��=��ö��6�(#q��Ŧ۳�Ɯ��ᕱ�}�	���4$x�R>[�6
E#�|�w�H�R�u=̲*�3j4��a��>�|�$��lvQ���0:�@�M�ϔ��b�e͊l�֌��"l�IW��V��/�7�,DD�'��}���ϜT�k�b¥0�D�A�(��A��e3EuU-�%uУ�?���H�J��H�rX4�sZQ�(��m�D�\!�=��C�G��ꋆ�� ��H�c��p!n��f��-b�bQ���؋ǋa��ߣ5)d�Z�7Q�z8����t�*M�|�Y1`�Ǥ>�|n}�,nnǀ�^hY��h�X�HU��WU,�����"[4�|��OF��� �����R\�t��i��1�`�c~�,�)�2�|�B�&�P�! H_��%'��㎎��iI ���L�U�L��uP�%8��әK��7�LXlI�?+�t��zv\�L���f]Ǟ�B��g��ڷ�$���<�A	u����l��{��A���� ��mDt�K�|#� S~��6��$KE�	�L��%]��Ra������ޞAX�`�6�bǝw����0;X�`��'�F*)�Q�����t�k���. WFW�� ���u����n-eI&�k����r���'�0�Z�ԆY������^=q�1G����@8^hÒ��5�G2Z@�o��٣c/��(��#F��xOdKI|1n�<	-�f$���������K�!�Q �Hզ��V�������=� �4�d�z��"U��d�C��G>����q�K/�1S@CMo,X� A,�h2@��|ɠ��ȡ�6)Wys����Y��-�J"��$)�D$h�*١X�LaE H�g�"��Tr��tlNx�:�E�����@�lS�"8x���#��1|���^���f>ٰ6 9}V �}�Ii�78I�E	Ѻa�[o�m�#uM%�܎��JX�F��f�=0hض(ī�s��{��A�A8D*��Ի��{o���C�TD!�6&�.R����PʛdUcq	�	l�Ŗ5f4���s����'v��|�F1V�JS��,	��P�Ed,O^&\	�����lwY��}"�췒i/���~��ğ��8wR�c���4&L.�6�:���%�ƀ~8��г�B�b+Z�A�e!⥬1������0̣�h,�S
jM�F�~��C.Z�s�b򔻱�y1��q��gMPR`̲ix�� D)(!oi��tc��>m9$��PM�:,!��S���P�GQ����x�g硵��d=7��\�R�����L{�@cƬO0�� �"$�e�E�i�I��h��?���xb�2��td�<.����c�]���`0=�%���RkQ��x겼F��S��xV�"�&`�$XW:_�=�`��tA����w�I7"t�^�9bz��kT%Sv��=�gϺ�&YK��JƐ�ŰU����2��8���=_���{�m�Y�m?3���G�rS�q�ؒ-۸C�B	�I @�!���mll�d�@(!(�dzI���EN�Ќn�V���g�������[�7�JG���^K:��=3{�-�{?�S�(�jT���$Km0j��;�i���[�����)�T�6��[��p�H��Y�Ѧ�����g�b]r���P4^i��h)��D��d��[�uB�u���2�� ��2��Xnx�b@��k�yӲFG������i�*�:�vڭ�W��s֟e�}=[�	��Qk�LYbL��U�ȲV�*�)���s��Q�������f^�<�ݣcv۷o�Fc�z��g��LN9[ъ�J#�f�Yg���bv�،��Wm�=�b�i���k[�8�Vֲ�8��Z���������3h�S-�F����6�w����A��G[Pl	�n#�G@��U�d�3'�z@C��rm9�4��A?�Ctar#t����hRć�#�ع&Z,q�8��Jb`�S ��B�)E:�9F;8������(L�}Ӗ�V��`'���g�� ?0�,0a��jZ��n3I���m�IgYr��7�1��-+l��JT5k�����'-{�v���oي<�z�9�U䈢�*�~@�RK: \���䣟d���lk6ˆ�d'���|���W�򕞶���G:0񼴷�a�ݖY7��!_Ch�u����1Wh���/��l��B�|0WB���8�p�Y��n��5�-�Yy�~kc�Y�6�Y���L��t�1*'�3Nw]V,��-'\Ӱ�����3]��ZM�R��d �d�֎�Z1!�����۱3��܊�=�vD�� Hcڦ�Bt�U��HR��+�?{�:�o����,�;8;�-b{ۭ���N���;�� D��Г,Sق(�Pk`
���h���*�H:3��}J(@b ��������
`ܔ+�a���(��)����a�Jq3���M�B�V�ݚ0���=�^��ㅯ!�o�z!=7��g���C�����$ɭ�6����R�X}��x��O:�F+��N��.�D@Q�(m[�N�l¢��nw~�VYfլe��3a䈘�R���zo�j��ѶV#��Zݝ�ĭ���XgUl�pᢧ�(����i;���B�*ڡpt�cN�7[�/6��~.�\���^���΄	Q[�}��_d���*hmIl��?�f�Ǌ��Da�y�H�(v�H�R-�E�7��DY�'����L�u3��jQ�|��#�05<|$|�����XEX��]vb��Y�=y來��l7��6�YEC�]S�Z���^9l��%vOOb�굶s|����h6�T��λ��{���#�p<@IX ��*��2ay�(̯�7��	��pi�������*��sТU�[�\�ܫ��Z(X8�)�DV2!ll�%�P����c�=�x�M�h+ŢsM�?2Lx� $wռ����m�1e�(�f޲��^Kk6�w����*ǜbc�A�`���|D����ylڶ�ل%?�7���;�*ʭ�6�ؔ�@��U�"�u��Z�8��k7���h�V�pPJ꡽�H>�l�E�Z�X��������ąLx6P�n���ƈ�,#c�s��m�4�r&�_��w&��*M�1�8H �JR-k����{�e��A���L���DE��Jkd�W ���L�[9[掙��s^l$
S�xm�E=l��;)��I#��rb��Yê��f&XےV��%�Ț�������M�׬���S^��E�Iu0�T���������1v����Ģ>�X&�H)��b�ۉj"t�AP;���0����~Z�q �$�0^U��>�~Ђq��P�ó�F�@E�1E^���LZ (|�@ AX��3�p��IN`�y�驤XSN�p(�~�?�Y~���
�iN�L�p�n���F���;��;�b@8�f�j�[W�9�@)��M;,����̏�k+Y��/�ʢ(6v�a�FMw�E�;D K��$�Z��l,����Z	�G8�e���(Е�p  <���3�X�@k܆��{A*A���|�;ߴ~���K����}��lot�����=zzk�6C�Ll��aI5�v���bbk2���H0A�x�Ҥ�t:�I���8K����7e 1��/ ��F��bma,�B�Q�g����N�%xiB�Q������#�2��ʽ����,.7 �m�V���p��y .�//�<�xFb�7���qd�8��$���#v�Lj�b����641i�ֲUa�7�'�nq���m]�Ҿ>��ݽUk�$����ε������w�i���@'��{r	��")�[��_K�l�?l��
�(YCq���tb")���&�⌹&�Z��(B_J�XA�@k��8�c��rM ��"3���9' V�c�.����yV:9��]�Ŝ��z��"���r��s: <>1j	�0��hV�]�j;��-;���[#!�0r���"����#�~�&���3ូe��I�Va������=:ك�� B�<=ȭ���hi�b�J��M�҂$�J'�g���CR\C����!g>�J��`J�	�G����u�	VI�48�8�q�g����3g$_��$�ʢ(���W_��e��󪧮ڽsc}rt�(;k��d�U��i���� �9kPiL�T��=��T:���PcQ��������I�p���|抛�(�,Ei�����\��+C�<.0-�u0�D^����ck�2S	05�`_��L,C;�K������+>i�+^]�ZϮ���ɦ������)[1=i})Y�5K���"P뵑�j[�ٿ��vgod��56�hYk
�m���A��������1��O��b�J &}�s���9C_P�A@XrD��uX'ז<!ǜ��ø���}#9���o��J�a�B
��@Mǜ����M9���&�x��yf��*�IG�� |��g��������y��Ƭ�vTV�aϾ��Gg�!�b�UXЋ�9���r��|��;�a�w�����YA�R��m�3_�԰�,C+d��� S��?~�l�+Q�#�t�<�,|���|�����2q 2.�����bb���"s�EZ a�2<��5TIN�͵��+�w��qM�cT�L� PO�37�|�O>��=Ky�y������ؽe㊬qN��0vֈ��5��&�њ���!;�<`g�X7!���r?���`N��w�k���^��luM]O�Nb;4��ϺW�����S������ߙ�Ej(N�"5����e��bLg��'~��LlX	&3�h�L-A���Ľ�!Qɬe6\1��kϜl؉��Sǧluc��r���qݲ4�
��R����=X��=�5KW���f��F�z*U��11:fqT�;����n�>icͻ԰e�#0py���{��/�jCK��`<�s��ń2�=d�jG}�~���u
�	b� �r�s�	k�Q<2 ��&��Zs�ZLx)Z�Ϊ眹��䞞>K�G4��k��7�m�ն��Z�l�>h≉� B�*x[Lzs�ik�qK������_�a�+B    IDAT:ά�Lx���.�
��y�c�ѕ�(�q���\"�]�2���L�tiG�!]Gc8�e����g��RҖ�<�'��3���G��0Bf#�r��ƪ+�xU�6,��kHW"��-�c� ��`�9�.Ϫ�'�_Z��o-+��Ʒ<}�ևoYg�4[3��*mt��ƛ�6�r�w�8��}��	D�p��aC�J(�W�dV0������En>��shl�I��ƕ'�c�NM8�����:&�âZ���2��yf5�s-�w�Ee�����8�/@�-k��������<�j�bY��n6�Iw@�՛X�J��C1j�6�vB���	[9M_��Yw�fy�I�j���j�eՐ}�?���m�g��pD��(���^�!;K#��]w�=�����!��Ć���;��X`X�'lsZ:�"#�%-�0�r����s/��:�/9��o�y��&�D�$��!˓#�+:Bm��<����WY:�p�U+�r�M�ŝ��l��$���yVԥ��=QݶWW��g�o���6�5��}�0�p��r&����6v׷mMlVO�	�V�p��I�ZRK<��,I��9B�/fZ��j8�$H,�I����T���F�2��!��31z��1NȘ�KV�|f,���
��(8¸;t,Ϣ�x��1a�; ��8�.�A���1w�7��ۧ�z��B�~>/�Wmߺq�=s6�%Ӫ)�vf���ο�v��s<�3�"N:_� �י�Hc0�y��MHb8:^�N ��_�r_� 0�I�ɤB��%��ΗY�Ux�FaPc��i� �@z��ib|��ꕒ�Y��u ` 0�zp��9���{ՙ�0/t0IRL!�D=P���P�E�q�Z�e���(�ά��6����q��N�b;zt�V����ܹ7��"u��V�j#q����G��p����nzl)1�+�\~ ����羻|��.3�A�5�e�p�$=�A�R&�,�V�VR���h�0i~�@!�HÄ�@Ӷ���9�c! sK�~�P�8TB	Yk��X�@DdA�SCLXKOq�L`b��)��n�f�Ln����B�Z�z�e͆ō�����ڨUmGm��~�y�>�D��;�x����<ށZH������6qwᘫ�g<:u)��@f#���d��#3>oD���n���]�նZ��8u��\%iHㆶ
��5O��c��}�o_��/~���\���}�+_��~����N�*���T����¤.R�T$���*�B�,�|��jn�xd���7�p��.+?��o�ڑG6V���'���i�0L��S��_~�m|t���>/����>���19�ƈ��Y��>`U�+�6(c/zы�)��G��e�]�E]�������*3J%�h4�<��I^�:#�2׿�,*?�9l�� ���֜�4K�V�&�jN�X��
Ḻϕ܁עj'�|�#�^�Ɏ�[���n�z�)�@A�Z�;J(��<@��8��Jl��{�Ln��96i�hR|���fI'�8��Zݶ��m�����F��A�k�SO_�;����B���N�Lfm��b���e *���{���߀%�(*|M�H *G�E�����9��9��7,,-Қ�_�V&�駟�u�x|�,&l��(�M ��ϸw@�	��Z���!'�8�:���d��C�Y�6rWR$k G��i�*��k5��-����xT��a[s�k��X��P��RƓWHB��2[�OYv���]�)@8���̤3�F;wn7��q*�t�Z�f��Z�W�#���!�VO[sjW����_���ojk��f����ox�k� -5G Vj���L����m޼�ﻛ ҟl��6i�3@��f�ݒ��?�	x^���Y�X�p�e��n��e�5����[��
��v�QG���?r���w��o-��{;,��W?5�UޏI�C���(���(]��X�^���yN;�E4>�b&�����B���U0�7�Zq�p�6B�2�bxp��^�[�j��֌բ�Fwo�tf�z��5S�	(N��׏�#��_�j�U{V�>s�nY\�ѱ	V�zO�)�ӍbK���8d�,��
�+�<ڵ۞2cvR�׎�lZ}|�b�����H4-gq���ց��f2������Bz{|_;j�o������% ���X��i����l8F82���Ԏ��+��\e�J_�0�BU��b.���{ca��6kr��z�#��Jh�,�b9>a���l �ǜ�qó;#$��i�B�pʚyX�ӟq��F�аM�O�Ӭ(�Z�I�؞dȎ:�\��z�M��m
*��E�G�,JS�6m�w�n{��^'� \DG����r멱04,�&V���i��}���<��x6��H��L��]N�l�7~�7|�-��E�J@ZEj�[,��_z�.�^1�A�w�ĩ�'`c��������Y0CkJV��Kƍ�+�2�@̳R���"�Jy�EѦ���=oYv^���[VX�l�S��s�s�=�%��w��_���Y���		�0��L+���xp@g
��AC2�1���a�����}��C��9��h����Š��`>��a�l�]z��G���/�'���&���q�͌�X_5���������C�En��cK�VZ�w��9�ҨϲJ�mٺ��vl��`ș�4�d� �}a@ވ�	��;fϬ���k���������ӹ��"���Jl�(��������^m;v�q�kR;��f�w//L�'֣	"�U�}'���[d�hb��É&&$`���'��	�д-�v�0�K��5fd��J�P�eq]�h!���a|1>���&���Ҹ!I�()|d^����p�96^�hj�8��{��W�cםg���)���L�2�"�-�2�[v�7��v��CF�JɄ��[����'���S�̼��I��r���g{�lUʣ�� J �:�SI��A������O(,���bA�ve�/��kQ`�,���2!�n�G�w��#����y�+�����uñ/i�-��<��[n�ſ;��Zqo��޺� �&�r�#W歳(̀���+m`u�}�;���W��a��d����Lh|4���Я�6��)��P��.�*�'�U��?�4���ц��|zp̙��:�T�V%޹�Y++6���^i�}��OY_���b���ZV#<��"��`E�,i�YT�V�g���6t�S�	�}�m�۴i�kp}�U?�A�>��ĥ�I8{ r#ʭ��cy�i�Ql�񫯲��,I3�խ�h�C��FaS��Ib?ٺ�>�7_�Q�SkuOÆ�T������r�䢋��O����ov�e�+>@S&?�$&JOz˖�v�Z5!�N�<���Pp=��U_jr�R�0��~ ���|.0��%	�����31D{hR
�%o�����H��zv�AD�_��0{�|��S�*���l�ն.��N9�,�)� �@�"k٪,��އ�����o��ﱆR�0�"�O��S�b�؉	vN<�?��Y������7�f.���~�ɳ�|��ޞ�J�ô/ɋ7ݏ@=��5��7J�^y�΀a���W� _|����Ӯ3|���4��}��?A�+-6�2��"b9���X�`��?g�@�Y�J*�[n|���� L��ac[7�&F�A�t�;�^��+m��#��;~�����(:����3(L7U�X��ѐ8�ІE�FD�{��^��0� ����]t�ׇ����+71�@b&ZqC����o�Z'�b���H���׾�56�_��9a�q�vo�w[o԰zJ�Vj-*�Q!")UL�v\���[uh��}�5}��^{x�N���M���E,1��AQ��zl�G��qbc���]��W�ꕫ��V�p_m�\�E�-����s���s_��MLO���a��ٕ!q�6��"��9���?�R�ir1�Y@5�Hb�$��N���`�i	`��@��� �P؟�����LL@���/�R��f�x���*$�iBr�7�����P�ǽh�`�`�!��E@4S�5�,��Tg�����}bi��.���l��ô�
Ql��X�S�ǿ������bl�n���.��-X|faYF\w!�M8&^�s�C��������r) �͸a�9�?2�{ �ō>`<�7�^��=��p���M>%�@�s�0�9xE8.��x�,li!4�j喛��ۖ�׌nEv&c�Y�<�^���m߻�v�O��-�='��	;
C�ԑ|���ʢ�����'?�4�������C����װ㗼�%�z�������WZ�
�I� �k_w���,jOZ_Դ�[���3�,oY���WN����.�78�i֎�����m㭛mz.kΖ �a�Ԟ-ct�I�{ѡQ��e/��׮-*��5o�^ �ÌjUkf�=�Ӈ���w�w|�������0��OHL@&b�F���߀_ ,p-ڭH�`p�4%��Ľ�ó^��	�Ra.��0����ώ]+�HzF]G��k3I s�0�j�r4�Pa�R�`�O���-a#���cR}�A�>i�ܷ&9@����������j��6�(,��Ͽ��F��`X����	5qa*;[����}�KvםŶS|�K!!x��$��\ �yC�Qʲ[�AX}�O1ae>���L�s���H�ā�ik�,������Ɲ�7c#S�`���i�a<�	��5|�w3oX�q�M�ZZ�$���׽{y�0s�[޴*J�z�}v�ΰ�/��~t������Z��0/V,4��ix
@�B+6�0 h:�������h<4�0e�yp&:�R�Ť�o
KÀ<ڠ�-��R��e��j'�NF;0�g���W��@ݬ1a}����齖M���j��r�mO)�=��Mm�aFT��/v[>�ֈ������#�3�.G(O$�lM����	�31�/8�<[�r�O�Z\+��)Mo�x5Ҷm۹�n���695U��E������	�~'�|��4O7(3��7���a��'&$읶���/Vǳq-�$\[{d�v����=�هLD�Tߊ� ��������sM�	��XV���Ua���!2�CV��@ L��D���}�z�^CB �~�m�u*���*#�������I�:ŭ
^$���ʨ�<���۾ioy���2�C�`6f�O1aL�n�%��d.�{@��B9��º�����M>!��,�ZHO�Ї܊�8=;�#9��4Db��z����g�a�ϸg�k����/
�ݺ}���fd��w����6,_��#�<�ЦU�n�iLu@��+.�0��V`1at~W�Q8x�O|��	 k�Ya	�E`R���/v�ba1���\@��]8K�9�8����u���V�,jLXo���	WҦ�F�+��<59��F��_���Ҹ�ޱ�6}�3%Sͪ��@��͂	�l���SE�U+�}�+
Lګ�� �9,j�T
5���ωC�V�l=�pk��*q��Ԏ\SN�d����3�8Ma�:`T&c��,_z):.\��59��2F�L��Ư��1�c���Ɛ@T��1S����!��$�;iC�_1M}�x�Ox_YWb��a|b��O	-D��g��j��	Ÿ2&t�.��-��νV��-C�_	w[V�H���ń�����aڌ���:Y�a�� �d\ >K�v�%k��
4��|�!t|���j/@�fQ�V|/�@���c�nYv>��p�ѣ�l���l ��pʱ'��_�2�#��.�?ǔ�I��!�#@�ae�sF�&���ԧ>�lW&.ǱZ��ot�x��������W���>A?򑏸�,P�х �s9�y��)X�<4�o�{�ڪ�ׄ{��3a4as��Äٷ���គ�c.��n����mőO��#;v��[?�ż)��p�	�Lt��� �Yy�Y�t~�@���s\j�r^4�g\s�]p�|�l9�rϚ�j��ݤ���`j�#�qM�E}*kF�mh���� �q�Z�E
�C���|��o�/���5���u���$����p����I�P��2?�ǋ���g�M]HZ�
��X�0�Xp��pұ�R"U��+3]V���@x�L�@@X}���0a����|��@D% �<#�'�g8�y�(EhgA�|<�5\�4� 9c69B�E�!�q��!�@(G�yފ���_w�ۗU����wl����+��1k�d�yͫ��[�{?�ow̱Zs�au�&��V"����F 5zaj����@f%�-˩�b���qڠ��Z�tP>+�+��a��q���Wmh��)뭴lǖ�,)@��o�ʆ�"��� 4r� �n=��Ӭ���D�u��u�glz� 5��o8��{ͤSYɒ��{�ܑ操h�>~�E���K'���U��W�(4dXb���sorӳ0����Ҁ;�rɆ�������^}�1��NOw�:�Ȕ���p�$	z-�2C��!h3f����P:�:z6@͙f�8$���P���"8� ѢP��]G���i�Lu"��!)��j�7�T���(U4bҘ���q�X��E;������4a->r��Mń���&y?�#�����4a-���M=����N�ue�9�܀#֢ȹC�~%>WʱH
 ��S�� i���p� �D��=�E�d�j�z˲���+޲y���%D��=C��W��z�k�����5�a�@�ۈF��Qd:��P��TMڏwS��u�Nۮ5��q<l�kʘ�M@ŵ�4[r��pֲ��~{��^cCu���V�R�������Z-J���A#1�%�=�Ȟ�,�)�^���a�ꈧZ�j�Zݶ���L� �g�h�ζJ��:@�v"�j[S��平&K�X�5Q	.c��}�q1MڃDwv� �C"C;�m!���dR��@N]�),g��_��~
� B�T��7�K'��hu�"#6%G��s����X��� 8�F�PH�>K��؇7��ߴ�X��D@���;�̘�Á^�<"����zO����e5�m	������3��� X�c.4�Ŧ�A����|�#ǜ@X�,
]{� ��[__gh�n�ǰ/%)��V������lN.�u����P��~�2qÅ����>��4M�7�x�[���O���C�����t 4�f�yϻ�.�������'k���e�,/nN�U7@� 4���̀&��<MT~�L���|Ql�L��W���Nȑ:[����V���?蓂���<�.��|{�S��;ئ�I�ڻ�c7L�R�<|�)\���Fq͒Z�E�~[uؓ��/{��s��w�u��~�h��v�ffx�a@T��$|��#T�M �-)����ZB�u2���\���y�P:'dܳ�е:��s��_��^/��K�!����Z����Y��X�B��sHz��bބ㑬:K�`�ra^J:�3@�^�x�����U�_h�.�M
g�B$��H�S"��o@����c �*�\��9�ƊC�6`�UeG�\IE�0E���A��_�Ӑߡ,�馛n�j�Ax�O7�Ό#GD��TQ;��g�%�t��{����;;���sS�):A+4��F6��j�@k�db<�[���T��*���H����>����B ��Ť݉�ʊ]*�w<I����nN[N	 1kY�R8S�{.�+�����Ψ��Z;K�V�əF�h�P����1E=� �uO�0���J�G.y���o���ŒP�����<��7N��~ ��|-|�\�o#��ZES.����4�	���_$:��%�%q��x���g�TVQ!��3��z��\t�ԅ�d_�H��/D551}q�N��L1S�E�EDa��3�2)e=��+W�k�cX�<#�O.T֕�E�7�����e-�^�w�����s��{�����U����֝b�^~�mߺ����d�bt;*$�����y���`�$|�< �)�H���f(z��>�1�
�g�h5J�����&���)_���l�AW~�`    IDAT�d����j������JU����b��)Oi��B�����1�Ez�I͊�d�N4ݟ����췀S����r~��&�;�ׇ��������Z~��@�쁞?_�?>+,����H����^���C e�IǗ�S@�q�����G��F-0���_j�b��f�V� �A��3��y�	��_��_v���)A�$~!�D��z�~$e*� قci^�K8���H!�'B��k���S�_�� ·�����ea��_�{��3��R� M8����	§�r����}���ǃ�)�W�It,l��A��8�b`��e����ωF���O�,2������ � (�=��P9w:�
��^Zi��%[8QO�}�<5�C�e�d�:�_�}���iR g� �׃vH�E����g��dL����u�`;b:� �{|vG�(�н�K a�L����?t��h���<�s���s��/����|����)��s5�B��W��.�[> �:�^�+�� E�=
�7rȨ%;Y��U|HDE��983'e�s����j����M%9���sN�#����i'ji!LӂT�1w�5�\�;g�yfQ�j��y�	;��~�P{fC�5ת=.GP_��5�~�Q���s�SN�`����U$��A��4
� N
'��F�q��ly�a�46���פ���~�������=��"��wz��4
����=e�I��*kC{s�����Yg��"[V[����)}0��m�`�Ԙ��n�b����� \<�����QW �>&�;&٣��r�	;_݈E��C��X�a怀Q��T�m�C�C�P�_�'s��v�ii�w��4����&���,���Y0V�b?���|���T� �H�BG� ϊ�8cpGa�r�GH�X�+"4��p���:�)�~P@x�����ҙeI���@��Ɔeնo8<��AX���(L�7�,K����1JĔ�C�`�rX����Z�ل�:�94���C������i�-d��oy�T�V��L3��)w�%X+��v �b�{^x�=�+���
zSP��3 �`,>��q�k=tt2i��7T��ھ. `>J��ޢ�K()�ό������<O����y���@X��,kS�$cO&{�a���V�I|̓Ї�9�<�$�9;[�-L����-���:\,n�Lt^x�����l->
���/JI��K ��C)�R���s�vl���t�<��O��]���eg����4М:�ZK��L����#���# �f��:�02�r��� ��G���W�)�Rv��,�.	 �zj�)�� �`�P�J@)�X��\��xY��öju׆�S�ʫP�����͢�O���J�I��;�*k(��������-��d('�&��i'C�ܩYϠ�JY:KgW�y����`0����"x0�m�k��[���~�Y�k��֣#gB�f��s�CPS"�%�N���;�$tg�q�:��clUa���w�+ic!'�AH��W_�q *�P�x�F����|� ý��k.�� ��Y`�V(�
CS vpK�=�Vj��<��������:�n�kL<7���w�(k6����^kΰ�4���*�m�i:��������H���@�@N=u�_ܯ)yL9&�]ך��\۵ȣ<`-�+O�(Aد�2��������F��)���:c`�e/!YDphq�-h\�-�/�z6քS�5��ɚ���kM�\k�I�x�n��~ޅ@b��Y~���х�ʅw��ShZ7!q?F�-T/�c���V��\Q��0T�g%��:�LXm�X�:�[ S�B1�Pn��h�\.�2,�S�V�d����"<�,�k��J��x��#��d"��)�
���kkY�������5;�nn�<9B�y1�=��|p_��lN@��Z!�٭�vj�e� u\��l:�R��_;OMݹ�N�n�u�ɱ�{�u��E�t���@��������r����5�">��н`jᙏHB	�ٚ�\��	�J9����hC��)� Kh����Gֵ�g;t�8��n�� ԭ�@�����T�� ̖��\s͛��	�����z�C���3�/Ą���k�-t�RL�C�Pj�'V�5�Ckx.��^;�����>Gy�X&\�T>{��W�� ����ڍ��U�L:��"���֥�n�^��r�C�j�C-��jEO��s���BdO�5�nv<_��:I��]{�o:�3v.����?����U��mj�\81���\�B��9���>t̡8�O�Av!@},�.�J��k���7� \*���U$���5��n��bq!yb1�8t̡8�O��Ɠ�������#� ����Aᕻ��2�:����l���2�����x\��C�j�C-���c)g.Ĥg#��ß;�r�� <��vk-!�.���5�!Mx)C�б�Z������n�Z�.�Z�Ơŀ}x�0C7I��_{�o\V9�舵;��35vA�'TMLZԂ�X3���D���d��nN�<�VP��UP�c�����	���-�U%I�|�z��}��Đ'�P\���L�ӱ9�%jf���ۻ�W�����Sx�f��y�����w�p�({��4�J;����u]�s���m�v;���<݁F/i�+����Z܇>���ؗ�Z$�����X��<%�h�������V8ǦiJ��篹�7.ktsk~pc�����6����ay�0����w	h�:;'(B�1��<��=kH���X�Ұd�i�p���� �G��8O�ε�����jd�a������S�49B���Q���I��2E��$J�����!lS��HR�}j�nֱ��:�¸P�(G�����*�	STM���+m��?�P�z�i���3�ɭ�.k��'�ND��Ͼ��|Ӳ��\�cۦ��q�AiF���3���yl5�ޥ�Q���\@W�Ȁ$����	�_����Tǆ)�4�R�<�&F����C��Ɂ0���r63.�䳁����ͬT} �0�N-c���Rjm7�	t�b��\��Z���|L����3��c�2�4�*L�Vv,��wҭ��®�WY�*��(�X5�9�td!/��|�6����иA(�!���~�0{�� <q�EY�VD���KYR����P��njS.��ԏ��7LcQ���q_�ܥ���k�K��򷵚u�
���TUb����m.���}���w��!����R��{������)�R�J8�BY��e�،,�pﱥ����X��݄�6`Nt��`57���X�Z���2a6V��v<P&���*�V���9,F��z/Q�)T$i�e�$�Q;�RQ0��ƠԢ ����UyOڳ�:[�eY�$��馛޼������9f���[�ugsa/e	�5��&\Mjv�	'y�3�+�h�Q���:p�S)e,yHm����:�i�IA �F����W\��Qb�F���O�a�}�3X~Q�	'�lZ�B�;�.!�����􋙨2�Y�a23�AX ���,Qas��i=�PLU����'��)|ń�
�<,��f-��+sB�E0lc��B�R��\����s�����t[=(�h\h�ƾ�����,p��z�v䡶�dRmH�ߜ/��a�����K.q�e)i�7�|�o-+����{��-mN"��f�3�4m{���/�~�g�����������F�K=8�9پ���x0X�W+KI��^��Wzaw�
�u��h��?��?�5!l^TB�^l��"�ʂ�	�Xf,p R45��-�P��<��� �S�Zf����*D�E�� I�~�U�:;Gk�w��$�¶�%2�(��%�} ��Rd�g�x�>v�ئ��`��!�9q�I��/��S�}˖-N� �b�c�	
�����n�+�qmI����R�禛n��e�ön�4؜��eq��5�v�e�k��ēO����η�Gn�X; ̍�TXj��P����#O�` �V&�����~�zc�e���0c���a0����9�r<�
����O�	=׽w�2Q�Ye�a��	���4������K���^ĀB=����c�'�"+�;�B@���b��H��ؖ���v�0�  aɀn���l�k(��K�K�'�`�<'8"�J�jW9� i��9��]��0hD[i�����Gb� �oj�K,�v	¿�� |�o^���M���Rl�C�ZGv�i��/�ܲvn<��x���29U�Rab�00d�*�.+<��/~�M/��<�����њ�~ɁƋ�n�wgl7�=��-e��e-N�(*�jgb��ahW/�ζ�8���Ga䅊sk[�wo�7��"�p_1���bcQ�����W���Q�Z�F�� ����9�m�v3"iv2��eIKܩX?_�I��g�1t�! L��"�0��7�W��fN!��ga�Ȭ ����Q�I[�I��֡���6\��5{�o���k1��"a�C;�l`�!��De�7��,���� �]t�c��,���.�j�	8H��l��?��[c��ҡ�<o�q|��7�������9/� y>��ڵ��K_�[�z����?��[������&+�#�ѓ���D������V/�3Iit��Fg�O9���/������c����ڹ�^���l7,Kؠ(�8�,ɫS'9N,�k�N�V��_�E��/F��,�V��hP��;)�^l���Y��>�������J�e��[�1ױѴ�Z���zll�iQ��r�FjOY���le688�+8���B�Q&S���;��X� �U̖��3������|��*}�]R�F��u�O9>�n��\�(��Śb5�0��{-{��?V��BKAE�`xX~�0m.F�lS�������}!?	�ɑ��o 5��O�=�k�����~�U<����E�����pa]*s.;���u�s��8������}C����|�+�|����d�&�gc4 T_�9�[q��
sN>�dg����q=��q��c��o�j�A��m��	;W��k��֝e�{��ܽ���~���*6�,�]���[f+���I�1!Y��h�dx(�>�����4 �\���x�w��M��{��^�A 4�Y8:"��͞�YO�~B�z6�h�������f��a��Z�����e6lY�kI\3��i�a�5��a�Yb�%Va�O���l�;.ge�b����Gj'��am�f�eyϰ�6sKz��m��3V�V��L-����me�ϵ�a�X��ڛ�u���y��Ō$7	D���x�ٖ��arL46�\�������w�f��ª�������Ҕ!&��K.�ĉ�fѣ?'�����I���/�r�s.s�c�$,��ER���/Ӿ[c^�G[0v���7� �@���`�� ��	�8�GO�,#k�~9W�5I"�"��M�[`�ӱC�g?�Y�GinEQԊ�x�7���SO=ud����6��8��<�ЦYk{��f`�����?m��v�~Ӧ'g|�L^�'l�':�	��ɁHs�I'������}��a�	X���Vt�� bP�����X��Ă�[y�jQ��<��x��8q�L:I(l�Z֞�a��ڶ�/����G�bGyӲxڢ�U���ȗ��;9�EHiɄ�J�;�K�]�YT+wp�,NSk�UK����F4dI��%�j��Q{�I��'��| �PA�.E�ȡ!�L:$MS�R%�cذa�O\,��ǒ�<�����k��a�/"�"�gԜa�/�C&.��s�)M�A��4a���:�|ļ��gø�a��Q����a�.spbΪ��	�L 9N}"�N?�tw�}���������5�\�D?c�FB��� �Cb�8�5H m#�!��̡{�<�c�����]�& |�5׼���~��e�y�sS�3����f�x��m�5f߸�߭VA̮�ꊼ�nv�VEn�P2�:O��@`�������?��yq ��
�x=�Cg3�B��x���0{�r׮7�*���XiIT)w��,�&�'��<֞s�����tݢ�bI��X\mZ�'���w�d�	}cP�� �Q,X9{����\��l��&����V����rа�9�k�������oج�Y� Xd,�tJ@�6�G�,Ą������A{k��<y�e"��_�җ<tJ`�6 �r�).p�o~��@g�}�?; Ä5��k@�� uM�����jC9 ��cN��\r�ƽ��Z �|G�N��W��Ua2��|��׿��w�
�q��	'�`�_~yg�^���9���'�"�n���e�6����9����	(�T;��L𓍇_��W��iG�{L��5��`�sЀ5Ƙ[�c�e��������V�Z�Ե�^�{�
�a�p�^q>�����Ͽ��z��y��=c��o��v\�E�C�����n'��X��:�,w�}�_p@�e aJ��c�a�p [@����$Q�\�.�b�f��Ȧ�Ik�T���m��
���X%���l������c�lz�NK'
�7A��,�iY�`Ū�Ŷ���<~�[�ю����۶�ڝc҈ݛ娋͢�5�A�6�o���-�eo͒��f�8lV3��C���x~&m*�!dG�i���g�s�1�MXk)�MLv �2�9�Iʀ���w0Pq��9��#�}^���o�������	�L�߹��s~@X���Ó�1��&���#X��� E�m�{X�|�V�d9���-&�pB���SR	�ym�� 2t LX�ĵ�8�3�]v�[ь�?��?��(9N>(�	��/~�k��E�v΃ �lն�Ap��6�m�G`Hj��ԧlb���J��'�s��o_V9^�{Ǧ���s�� c���^l�}�y����۶<�S�Z���+��C�0aq ����!�����eT�kݺu��7���$�$���4 �Xߩ pX��l²Jd�z�=�����ZOo��m�Ѵ�c�p�����Ǝ�Vi�]�h5'-%���e}+�ĖEm�-�=��� ��P�x� a�$��u�2��5sL�Ul:^a3=O����f��Y;^m֬����Ծ�w_qYFN-|b�1a&&�����ĵCY)���B��cp"-�ޘ��������W��c]ˮ�5���������7��#cx� ,тL���1��$'�m��r�s�m�	�9b�!�s>}���w+����˄�L��/���}z��9c��b���+�饗:s_�YI�	$M���h���cq��8H#��c�>>�<o�qr����o۰aÞ�X[���>y��G64��E&*��u���_d���o�O~��U��E�1�r��蚼2_���,ei|��4�-���%F������J�ַ��l���R#�CL�*+W|��
p-�Y�ֶ,�,�*����v�ŗ���g-��m0�a���,�u�ٞ]MU,��Fl�hOZ�3c����-�"l� ��ٝ� a�+�S�*�-ɩ��g�����E=6��ht����Y���hX-��*�c�6����_g���X�&�b�0Z;�-�`��F�H�?�2���!ib��hh�qMm)�?�'V�&�R���X��Zlh'_����Br����Tp b.(K�$�D�Lr_h)Ѿ�'��C�"�\���C��9�(��a��ǜ��"�@�`�,��]���Iý �<�^��Q�;�ڗş�Xg�{���CF�P��p�m߹C�ҵ�(���k������]Kc��ʇ�l^i�s	�":��O����W�w���>K[ W⃆���$E�<�< Ecȁ�g���̅�i0���I�~�s��f��s_:�L	9����5
 ��v �����s
�)���9b��N�O�g���X2�ǲ1<f�j�5�զ�oUb����q�2L��H���V8�J�!�'{��t�&z�x�{l��j���#,<����md���zWZ�ƶm�öi�-�Js��2���N�ðhO��2@��(�+�n��̄�[̈́T�<��O}JP��d���?}�R@�c�J�pѓ����R�,�қ5OȒ��EVćc`��0����&/?O� }�3oC�l    IDAT|�j�p��a���_��_qf/�<c0&�a�������>5�Y�9+�Ϲ9�p>bi�=��},�x�y�Ґ,­۷�5�$i%�ʧ����߾�䓗�	�����գ[nퟙ<��nX_������Wٖ����A��乯PԐ�a���D&l�N�� ^:�ق�K���t:�@��y0)^���q���| �55�+�eI�</��9�γ�/�Ģ���̢�n��X��n����{���VV��U��5,�N��a5��Z֎�;��!I�j�p�� �e���{F�<�i"��L���DGZ:t�eC�ۤYd5��j;vm��}�c>xh7M"9xfs̩M�,&#�KE1����4�n��IqL(h҇�-�&� +[I�|6'�OZ�9�&r��������=�dԢ���#�����R����ʜV"�/�*�G��:�#s&�~+*�>Ww{� �w�Gڡ|:��=��7֏�p�6�关��q� �w������cz3DNl��E/z�;���	<P;s/$v�`c��"cY�q�ߐF�S�Y>g����_�ӟ��M�L�m�I�r����v�o����G��:�Μ�8�U}+�5�y��+���g�j4Z�P�xb�$�j���x0Y���á�`��������x�
N�����c�G3ؔ%#`�SsLK3��YVi9�ҺmX��.��R�)�Jjq{��{,�����Z6�����*�%V�v:cV���ê�ͨQ������ a_�<��@���C����fU��W�Ht����[{�6c��y�؎];PX,�����^����!:�1x?X �-������\d!���A,	-��_AցE�,��O A��<���m�8�o �v��x���с������~�/H z@�����':��G���x���G?��Ge�2��_���:I@� 7�����d	@�R�3�����I!�$�3Y��8N6�|�o]�d@xŎ��4��#�VWM{���8�t��o����5� ,�S���LQ�w��*i�����/ o�V8��I"a �)���/t3X�k� 7��!��{��k�P���t'-���ε�/��(Z�T2��^�w[4z��'�u&� �V���X;�*@xM͢����aq5�v	��Q�`����펼*���DByP�ØV���Z��K�i����Q�,J|�	�s�T�ik@�I:��B5���̈́+z�@�����2�q�2a`8|��$�[lsR����
��b�k�qA*��s ��b�1�áDԊ<�rl��cɄCfͽu3aƗ�Z�Ҧ��7��1�7n��G;]u�U��}���Xrh ���'���'|&'��QV���NEf���yqέ��Z�ǝ]N�8�6���w^��������j��;o�=�R�#�Fn�x����r��{k��ۿc{��u�T��<�FiHҠ��cN|�;���d^�9A#6��/��l����'��AJ�22�^ �=�q��(`^;����n�;�.-A8F1Ha»-�{��L�rĄYҮX-��c�%�yâZD?��@�9Ⱥ�� �Y+�!�c.+�
��ؒw�5�NV�H�p6�D�]{v;v��qhƲ�	�	��e�jA{����-
c��o��+�`EL�4j�έ��q  YʄY걡�p+�S�E���X�򗐀�sa��_���X�ɯ盭m�N?/9B�7�q� �u�n��O���6,�$0��?�tX+�p�X����q��״��44?���tb�C_@���/��R�7iǟ���w��noodsc�<@���e�{7<�l���n����L1xJ�`Ő�%�=7Xw�q^ד�)�ê"ݏ��Ӈ?�Y�t�M�'�h�l�'g _��>�B�T�%B��l(����S�f�����B��jn��a�#��,۽���أ#`�E%Nz� Ѱ
L8M]�)4�"Y�x�Cj0����d�I9��������׃ӡg�4 l5��9��>�яt������t>��оfa�c�	˯�s�Q��I$����d�md<���BR	��c	�|� J���XwH�[�O?��uc*S����Eb���ǚ	�ϸ�L������w�	kH�j�P��i+B\�z/�g�+	��"��t/�"p�9VQ"�M�0�JQRT9�r��]{���}��q��y���Q���P�jN3���U���/�c��ۻw�'+��t`~j��0����d��<���48C� F������Tx	�F�����A<���`Z��c��#�~~5�ن��y(�9@8j�#��{��=�-3���,A����6c+V�XқZ�Z�	�{Z2�C�ps����,f�T�פ��4�Y#^i{��>��Ԧ��1%�k�}���T�͹Js1a@9��	?� ̽�AĠ'.���������cG�C��c`���`�9�T��}|��G�3�I8�]8� a�5!�<�����_�LD%�������!��� bƳkLз|/Y� #sN�j�n k�L�B!���q"|�aI�\�q���u�D��Dj���y�F�����~k�Ax՞�n�Z�o�Y�*_�o�y��G�e�\nO}��;&<������(�a�_q�����XB�-��D�������;5�u�D�|�΄��S��>�U�2�(����b� �ǹE0�ֈ�,Ax`�f��[2n�kWc���ZeƆ��&��N����v�.�o=羞�QTS#"���URSw	WJM�hOk�LM��Շ>��t�9��҄CGR8�5��ßgt����,�)�i�L�C,1$
�0�1@VĠ���9� 	�Ysį��x.2�p��_p����/�Y]�7>X�9�[��$k��m�I{i�S,�p�=�UD6�X�)�X�)�_�D�(� ���H��e�b���gL%I�믿�ͧ�vZ�f��W.B���?3���6��!k����#���ϿЫ�T�&	Ńk�X�y`�[<�8�4�@�QQvV:�A�7�/`��8��C�r����}��sˑ����9b�q�!e0W�#.��b7�Jdyk�V$;�2r��>`�.�plQV�V%����:m+�L�A&L�Kg�D�)mY@[�����F%6�䊈	��	Q��m$:ڲAs'�t6XD]X�Μ}�`�s9$�c�b����v�-Ą�cN��B��h�D_�rR�����B�L=͇n=u!Ki��h���}bZ�З��u2��C�gZ$�Gat�Ƶȅ���d�z���&|�SV��WI�q��9a���r��>�`҄2L� Ua�*����5�/�o��^K�\ߛ$��������SNپ�q� ÄZS�Z�EloT�F���N��Xjδl��՝���Nx34�J#�aa-���.�ք'U�X��Z�X͘��A�j*�.!}�L8�T-w/<�#S�p�:���+<�"�T��{lE���?���,ߵ�*�5/{�&�5r�iZ�cվ��6eq�>w��Җ�+�sA��je��q\��OY��cʆlĞb6|���������d������G?�1DZ�d��jr�=4i�R���sK�q:<<f���Xf�&�)m��	� e*�1�m�p�R3��g�1ǘ����l8)�pqYʄY�cgc�ZS��-+�]�q��r̅���sR>�;��?m���e�"�[9k�gQ�V���\EbѶS�1�P{�f��o�qE��0[,&$Q�^�B �(�`�~`A��$�Y��9�ƊA��P�?n�⁤�J4g���r6h@i i ���x脜�/%L$��#�4�(���iIԴ���%�\ayT�(�ytĊ������F�|�KƫV�H�Ȭ�p�C�*}��(�S�"G[^��K[�E�(k\�#��&Q$8Sʒz*�3���3,>�Z}'8[Y�~ddrY@�I���c�Q�θO0 ���zʹ�@�u�j�Q	a�j�j�9M�p⨏%K�\_s,�� ����{����\�x�ɿ\�/'��_��x
�R���n܇�Q���e���A���b�b�ݖ ��/�
#���f9ڰ���-�p��И�Y��H��2�3����2���~�-��/��/����u�-���	�\c�2�wZI�h�������Ԑ���JիÀT!l��,J�Q�7��}V�����l�����c@���V&�,��c�}�l�N�Ɖ����0��,A�m�h�ab�Ҕyw��>\�1��uΫ�!�"��|���3,[>ѦmЬҶ<�ld�1a&��61dEcU�"\h{+����<�ؔ���K�FAh:s]9ESE�/���1�!�-3�X�/��J�S,5��D���̧��a�@�9����zDu&�8�� _��cT֡p!|v���/��4~��y�RP}�ꫯ~���)���d����<�4�pjUY�����%J�����>���2�H9v� lYW-&D-�a�L���"D-�A��ȧ-�4l�0�p� Wr��,�Ȏ+�E˨A�����Sт���F�ϩ���^{�e+N�f߉6� �~��ޑ�b¬����M�y'����j cn�?Ŵ���9� �|���2���=F�_�R�Z��.�*G�sD ��e��|�X��
L����+��\[	�}��jĜ�[���	/�8�!�MC��M��h,�3�|�mY�a�yI��tssi�����v����F�đ�NTCΦ	k%�3��.�@���>$I�˄�j�~h"9� �K/�ܓ!�J��ֈ��wX4r������[gUK) ��XTi� L�ܴ���R@�eׅzV�q&iCr��QA�cW\`�$ =Ͳ�S����0���yj���oM&�IF�$t2���>X�ژ��!kcV�_&��JJç_ m�C%� F�T(1i��g��Q�D���	/��1�YHHr^��#Nrڗ>�?#�x����A����1"���>d���"�K�-/dg;&���tȴ�H�� �CK�G�<z-(:����&_z�;����g���W"��	��6�&�Tc���� �!�sp���39��%GT]�hg0��ˊ�JdI9b�%#�Z������'2KҚeq�Y�� �#T�_���˗6��w6�$�W�k�gЩ��d���FO�lų��m� �,�ѽ{��f���^�2�F�T{j�G���)9�|E�p����`�&6!�h� �����7�^�0a?���>Iԑ�|���x�\�+���0a�@E�f tZ�	i�(���8"p��
�|���x��F��6n�ܦϥ�ӧH�:Sd��R���$-��]J_���l�fr�"fb�]-�"�)ZV[qLX$ܢMU0���f�{m�j?�Q��kU	�y��р�*�P�;�,11�Q���B :"�+%gv��뼞0�I%�>+���z��l�6�ɖUҊ��m�M�jᘫ�1iqMv[TM+��[��Ow�#.�Kf�;YSLq�&�a�c,_y������h��fY��Q@���̈́e�2Y����U���r�i��M�|���5�b�3i�Ì�WIH Oz��)r  `X8p�!�(*JYv;�y��(�N��@����!X`�B`����I�� QO�0���F3>�Ѩ���o�)���`GG,��"',V�~�n��cDFĞ�\Z��`�>�/_}�տ�sg��u5��թ[��i���!u�:�������D���`��SO��CmR�G�����.����]���c[,ݽ�l��!jq^5j-��=V#m9���kl Zh�*a��j�o���L�D̡^���m��\0e���h�'Z��X���Q�3��>����4X%�҃Bט�r|Jv�x&.Z;(8^+�ˎXv�Ez�yU��3R���1�n���:Ąa�%bQdn E��`� ���N�d�J^�| Y���IW�{J�R�������S���g���.�Wu;5�ĈC|���*`�v�q^����C��F�`�c���}q�u�V��&�LZ�S����aM g�e�p]S��YAè�j���|v ���m|z�*=��f�%qfg�;�֟��B���6PkXOk���wZ��Vk�|��vj=l5?M��*=��V�ޟ[�PԽ�l7.����
�}#ϝ+I�>���~��UkE+m�~���Zk՟b�jeв��G?���zM��[�_��~�U\���M:Ҡ�6���H�..���Ċò��$�����������c.�ﰟ�]
�׸�<~��)r!F�x�<dRr|jQ�I;�a����J7�}��-����B������=Q1�$%-���{~�%�cMDI�����g�kt��>�YdOq3ܛ�l�w�Eڂ�BB�=��Ӓ��x�oX�d���4Ԟq���nMb���g�S@��0Uוϙ�ܸ�e���A\#��al����X�a����^22'.��g�L����f$��@�������ZW�hU��b��"�!�	�[���ZwHXk�U�j���T��ֺ#n,!�(��v��������͏;s���0A�>�<�ν����y��|��}�{�ѓ�jé6<���+͟�gޞW���J�f�ғ?2�������4t�})�R����fͭ��Y�)U�2���Ŏ��O��;͍.a.�p��G�s�A�[ޏTSo�i`d��뻺ӷ~�5���z�>4+oo�?0��fW�wݞ��pΧn�b�A����ٌ�Dd��@ϧ�R����ar �5�/R>s@ǙT�d��B:K�C����&N��O�y�:���s1�`��1�J�@X������0�H��m� `��;֔���˾k�5LG]���0<�L<rue�jo
ޭ�8+�3 �A9�� |�����-����h���8k�O�B5�.� ��wDo
���W�s�_5�5���R�|�Bc5>!����T��I��q@`7�����Cs����ݝ���Ҳ�H�<|ߔ�ߛ��G<YB�!
����9]����b1Fa T�h��l�+q��k:X�\�J��4R�3m������Mw����4�wn���<��I�Q�� ����YC9n2�e����HhG���mTpqq�!m�̲��g2cLؕN���;qO����xV�F�q5�u,�8(f[��j��X����`A�v�(Q�6����x�5�hg�qħRg���{%�8��?JأP�K��w�H'���1w����Q&��'�y3�ޡ	+�\\P�a�N/bt�9�����gܪ�q����1A8�Sȫt��z-k��*}i�V�	�{�7�=u�t�K�z��<�r��Й�׺rv}v���~�#�d�����0[�0.rDd�ݨî��H��oY�(r���M��J��3+�5��`eϼ�ܬ��42ܕzq*��	��;��ul;D`G������y���'׍S:�����ц�e9��x�x?l�)5�F�|����e;D�}�m�q��� %��I�siyd��c�D;����+��}G ��y����Ĉ�v�s��&��vm��x���0ʛ�m0JL>�q���:����3����4ox�ɀ0�0;k�	Ä��p�O;�y���J��p1���r�Ƒ�ϲ G%��wݑۥ�+˶L� ~��s�B��,Fm���C�eO�>�����Z���	*Sw_ޝch�Z=/ި�i��)'ú&\�z�����	�yϏTEbIi`h0�V� y,�����ޑ�T�w��=�RmhG�&�N=�p��:C��� ,��ь�6|Ɏ�%�C���dJ���#(	XN!a�q#˩v��:_)I���"HH$�t:j�x#��b�`Tn�g@��8˱�c[ęQ��9�_���t�o�{�A][�;,'��4ͥr���qF�����ׯ?���,:�m݂&��2תEn�rr ��I��ȍ��J�NI�C�C��	�����F�GϽz�w�0�#�E��0�X�Z-��HwW��3�D���ONVv�����W��9�C��v�V�'��x+���H�N��ùJ��m    IDAT�r�E<p��Q�w�``뮧
@?RO}LS=�{G�}��4������ԗ�#�4<8��K}�l4�8��٥��LB���k�Q�ߨ;�3؟�E��i���kp�ZN�}6ʍ�ow��S5`m[���R81,�6�2M���(�U������	�n�1��o,�1�Y�`�-r�a�ܡ�R�Xvن<�P4%1��` g{5�0�I��� �c �V�����	FA���W�[����a��{��-7]6���ı@�o�G�$��RHC������O������
�����n�ǘ{�D�q�T5=�c�
��@h �f�uో\�Y�������Z����,��\�I�������`���2-'>���`��]����袌"�ew���ݬLN�Yը���]i�p�W�){�9���T�	�y9��3E�����4_s��؉4���O4����S:�:8���I|ﾲAX��Fg4�Eu�������v1����m�]��x Xx%)�7�x�V�C���f�Q��Ⱥc�&[�c1me�Y6:g�D��O����a N�û��㽭�Z�FR�O�]����not�)o|̂[}ټၣ��#�,MG�<O{`�,�t)0@L�#��,����H����F� ك�կ~uf�9²��_�%}����F�lC��:t\l0�����@�DO7aa���RO_5m��K�>��ޮB��W
�2�YlW^��f��sNI9�0����bۣ"�;�,3Lf�gw�kp�t���*��ix`8�)���]��h��3Ə�k QFh�c�'W�;DD�O��9U�N�DԣǺo�X˯3���d��8/- ���h)A"z�%b���l���9^�ԁz,`�H}4c�9?ړ��l��J�2�";��C`x�@\߈+���X2L���$�'F]���稍�GA�̎���3�}�­7_6����f���������@魥�G��z���ܹ{��}�ĎJ�!���cB� 8a���I@dtTSw�[������8 ����,6d�Ҙ��[��e 娅��JA���ʷ��b��w(ݦ ���FW�!d�P���G&��.'|gq�+��n�1�sfj`���8#V��oH��t�Ȍ�-��/�F8P�q�gnԈ� �0Y��y����q222R�V�W�^����������qo��eF�����>�ꛛ����%��}.�g�����<3Z ��;zEu鄃�`h2 7	?H�c�Q�6��F$������Pl�Ɉ��h��2��t|���f6S������j@)�߉�!18@�~&���0�S��3���v�Q��0��7�*gI�3GI$��N�Wv�t�pT��U��O�Y��� |���{���n�t�T[>8ԟ*�=iN����כ�?���'<6���?L7�pS~xG&
�X�W��2��T�ёyg��I�u��(lEr�gf����hv��yի^�+��@�0vT<��L�����=k �����/��>�����ӟ�tƒ�N;-�ڏ}�c�8i��'P�p�	YZ��%��o����p���*P�o�t_&<��U*��֬Y���2a@x��o�t��m˙2�T����ZZ�|Yz����n�rC����#�2Y�:#�9�@N [�8!��lO�6��xE��9�5�C�1B>�y��K:/���V��{�}��5S�����V5 ��߮]�6˖��H(Dn����gdݖ���o�L\b��g>��!���Ȑ�W�z��椁�q-�y3 PwvF�X�j���޹��9��d�	���+_yR���M_��������<t�=��fu9�0�0
�;R@�'��e:�ta� ����f$#/8�{���8H��V=��L����Y�k�o�ƍ9���?������s�T�d��ߌp@�$�j�9���~��8j���c�0��Db!��?��$����3�Wz���z}���s�ʋ.:�裏�c"�9��Fh���vå��+�g����:��?O��vk���'��0� -q�)����lt_""m[��]ՠ��b�w[#7�|]2��f�੠�,6.��d��D*v�ؙ����� }��~�Yge�ǌ�+_�J��t�Iy{�ؗ�����~p�햸; �n�`~#���J S@��	�u$�Fd�w�'�
}�=ц��ow1�p��犕o��G�a^t+ <�"�k�w�#Z�^�����~�����s�c3� � �a6�y�o��%nh��~�s�˕�s���>7ꄓ2�u�ע!�hB��͵�1�i�0s������	�N=���p�%�4��������H� "���,�e��A3k�M+k"}�S�p�br� �W\qE�>�ឞ��^|�9aC�fo�gEo_5uwU�҃O/|����?��t�/�z�}�
�ٳ�l�~�2@�QG����k�"F/�7�q%
�d���'���m�љy��)���vr/�s��㙹�L����k��f��0�8q�� ��_�H ]�3��
p� +�~�QGe�fd�=@��dʞK@ 8�}�o����+�+֯[wnGW̱Xc��o�l������R�қ���)�9�yv���+;���B~ (M�e��Z����<������+���Y��-�tR��Db�Y0�py'ͭ����L�&w��؀+4[�4�+O�r �剋����&w���fj`�5�bR'���$�����~&h��)�a�G� 4Y��~����Z��֍�pI7�s�x��g~��[2^�j���+6���Yf��n�l~}��=��'�bɲt�q�������0�,a m�/�1!F�&L��f5���e�\�E�`ʡW�� Yco���Lu�Nfq��IE�+��d���yqE���������@���g����]Q�#��������P15Z�hq��C� +�lGb{��h����a���+s_��/��8�8�.�i�;�w�i��V*�׬^s^g�#N;瀇ܺu��{�Ȋ���i�cN'��������?�M{Ι�����a��v|+���n�v������O~2��6c�,��F$e�mres'�s��
�h���I���,Nڽ�T����u�KY16�nq��<�{Ϝ;SS���J,0��MDF�Y��=&�r��/� 4�4\���0�p�o�;���D]�w�e��&������^A�V�t_�f՚s:
¤�|ح[7Ww�Є�ki���N:���Gw��7�=�Tzs�'t���&Y�s#���k|!�Þ��?�3�ۿ�[�B ��s��:(k8� F�1`׀.e� e�;�	�G��Bx>���j��:�����['N��aДGО�#vU��\�� ��^t�EY����?�#�d����?���o0�Q b��׾6�� ��nr�{��9���H$Տ�vf��)��ȘE��QЮuww]�~��7tT&����o��{��O�ф�Y��c��yp����t�w���"��K��� OY+� A��d��J�2�&¡�4�!`�nXhs�4䪫�ʂ��J���54f hW��PN��N��v���� >S�������������vjv�]Y0^�[VŲ�����l�1c�g�}v�	�����Fg�`;��&�� ��A	��s b���I�93(�b�.�Q��bnÆgw4�;�Ϳ��s��S�v�sC���_�����$n^�|���
Q(u�Ȯ���p<������ׄ�?�ъQ��/̕�bt^� �ד��f�\	CÙpyW3�VH���it��1���u&�{̲�5�z�_��;`\^54�	O��g��d�G 
o�۳�K�6������R�>��<�Ɩe�XDz��$n �a����q�]�'�;,��C̈́�%��G��q���wt{�%����o�_�JN-�F�J�?���)G�'�����~�n�qK�XP��S��0.� ��̱_#�3� \��9DE�(X�3�1�?'��	9do�����a��"G��-o,�I�mv���D��`���@t�KYC��e���L�`�Vlذ!K���Ӻ�;F��ۿ���س)���! ( 6�G��G紤���lj�#G
������>s����y��כ�=�,jh��g�K۶ݗ�~��t�I/O{�~��~��F!e�N	F�_�# ��K:K����_�r��-�y�a�/x�r���5k�Ne��LN<��� �o�FFD0�.ӦL�>��g���ەe�i�d�Tˍ ����͙����Uf��n(��L]���`R&'��7~��,`��'V�� 1��b�[臨�p.�{ Q��#����(�����ի�\�b��v����]�����7e9��-��3��N��f��K�����G�I}�~���0��.tH�V�e)!���qn�"�������z0Ss
��%q�X 6���#x�r:$y~�ɑ�ӌ�q0������kT��1F�-����5���
����=^Wϲﭞo"���xl9,��R��~��(�Y�гo䑳��F���{�R �v1f<ΞʳJ�#H��m�M"��%쬁4qd�da��^�)���8��� *)FGv�Z�z�ʕ� ��nټ��}�u�����#��?-YrDη�*5m5��Ί
�~K�(}�m7�V��^���F�wݷ��T������Z���t�TA�rǎZ�.Q'�Af���!vJG�<��&�',؄�+!ŭ���k��xJ����ࢮ6è[[����8��Ȩ_��ٞv����a�!�dL��nx�mI��6NV�QB�OJ�F�����$���	[X� ��.���?���!��f�h�h��F��.ᅷlټ���c���]��7¦��4��������ex yHqTعy�^m�(�Ȥb��=���P1�Л�q�2Io�6IT6��ow0���pd�J�*x���A�E0��z.l��L�S��1F��-��'	S:;*���L$�re3Ze�����|Yg?��>��ːe_q`��9 ��Vl�����,��
�'���q�v�ߝ��g��]�������h6�C��|����E��o��	Q[x�-���C*���Hv�U*�y{��jW�>��R��E?!�������Kv+iTP��9��ў�q�^+�����Kc廨�L��L�}��F�)�O��m_|n;��c,c�0{����k�S+CZ�aꋲ.�tNɇ6a��3Jmۖ���3r��V'����2U�Ҏ_f��]<�w#����A�ߔ�l/�]�����S��о֭����)H&�G��ܡ3�BWRg{Q�Q��l>�jժ3:�	��޼i�4�CԈ���P��+�y�{k�l���
��x��70�w
^��G�|���]��q^�{E��4��=;�Qv�^\�5c�.q�ȭC�7"�����ĥ�tv��#�N�G:A�rQkC�f���#{��Ap:۾�{��r�38I����?���U�5/�}N-Y�ٶ�ɸ��rRԊ��(��ygJ�_�g��c�?S�֫�R��D2��,�D$���J��yΎ��[6�ڞ�p��I�ၴ=��k��OIc�Ԝ�8*;hQ�N�Ai�\S/��0��זEG`�#�*ǎ�N�@�B.�� �p3:��Og�dY�I&�(�jL��п�y������~G��҉��`��N�M�{J:t�Z��$5��Q7XW��������՚�f5�2�*)	��a����˱�M��Hg�;�	��y�������@x��n!w�15�UO��	���L8�q����O�n��4����5Em3o��:�h���ָ��8�
�ց�6�8pJ���{ �a��>��G��� ��.f�����	�'L ��� z���Q����v�{�ʜ�҇�oY�ˀ mI�	��� Sf�T�s��>��������Y�ǎ\�GR�wfBq�Jh)�%�ҁywg0�팜:�e�\g�b�����,������R���U�N�a�ڞ�ێ��Ɏ9�-��	�h��6,&��,I#��� !�Ƒ:N)��N:�1�?Fi����S��`t*HG"� ̋�ynS|�8�!lQ9��Y6��g=+k��I%�&uFAX=��pʱ��N$�)��κ0�[��e�W2 J���?=�����G�đJh&Z%[��,D`�5�g�����Z��c���S��T��0��ݩ#R�������X��uhc���|NyIሳJIbw�g�$1���sٯ��R������Z�~n�ʕ���7�ߐ#p�EM�|�lo4�+�k��>t�si�udgN�v�!��=Ǻ� [�3Q$n���;K��q�-��]�/����A\ո(&L�PLØ�u �h�>#I���eS�9"o�z�U�]7��8c�{�'rvz���������%3b��SN������75�K�_���e��o~s[^d#�"	�7� 6��~X��C�^p���X*�c�2��h��I'�@rg��g<�`Vf���vlD"!��>�6���[��OG��U0�@�ddƞ�3�,����V�^=} �(:�*v�8-K�h�3���\�� 0�����j����@
`	[24�����v��rm3�3	�x)FX��&d��> �&�S�k�0a�2jSiߩ���p~��|֡e��$a�h��?;ǰ��$A9L�A�#�Hc� [����`�.�k�\���xΣ=a��S�^�}h{ڗ�|�0�^�r�=ǐ��킢��l�ϱQ,��V}��~����ҁA����l6bV�Si�f��e����իW�:mL��
��-m���:[�L8���P��u���a�9�IX���z0 ������d(LU�6�9:*�ҹC;q䍨r�B�AnP^���7\[�w=�s�<e��� S��v����ߣגf�J��A� I�=�i���h����m~Е9����r-]~�3�%�����n�àMx"�Jy�=8�<����L���9���� 2�2�;x5g�o����,"�h�e�Fn�Kwww�A8�	�~��yC�O6:b,9����� qA�U#8����\!��P�*6B+&���Q^�̹���	�+�|yǠ	�1 c��YB�Ш�{����q a�q�kP�g̯@�W]	�DD����Sov���:�6�kE���I=�qw���EG��Xe���}۔��3 /�~�����3�5ϋ���V��
�9β웂0ύ�20�~?Q�PD[�n� �#����s<�Y�/�p3v@��rI�m�i���O���'�v�~q����oy ���*�,NכU\������@/w�����l��tZ-/?�n���~�ba6����Ɂ�@�5�N���AE9�c����܁t��=\�)@������O[I��TR��xw� �m���$�h�q���b���؆�q���oAK-U�Zߋ�t�ǁA��;�C��bߚ.K��-Gr6D��3;�)Y��r��>��������_|�i΢v����qæy��O���}F�q��fc5c�>���]��@��)_�ȷ*�n��ǁ��bGta�L��b4�XSFt?e@�Fa���D��q�n>˰"s��щ��g;gy���;�d������:���d�N�e�����`���]�F=��D�1��vv�qê<��8+⻸�7��LT0���#���a����P�Ѫ��V<>2kYh�-b��e��s�7�'~�Z�Hi�	��&|�ƍO�hRw6�\��f����@��M.�"D��м�HV���)T��+O#�M��݊I�j��{3@m��~�!�r5�������}���L�-�h�YM����0��b�ttbK��[Z�N�k��5T�G�=ֽ�S
�D@�H;�>�0m�2X�����]��\�/PF����w�j�\י�������ϙ��Ug0�%�����=Nn�k    IDAT�˃4��Y��"�Ł���@O=(��V��2�6�y�#&�Z�8j�J{�E$�M@x�T�6l8�� ���s�ϖ-�������Ã�T��Ô AB��s��E��e�cQ}��Z� ���S�����"��G��x�؋����	s0ؘ��%�t^�&E=��3�Y����&�-���=��*I����M�������E0�Q3L����zR���U�V�߸�	��d�q���UG�{��j��G�$c4���pu`y/��t�U@�r�dAXP4N�ε]`�w���l�W�tf�5�_�ڙE���c�g� Bd��PgQV��������������s���?��-�����"�����ܞ=ROO5�n���7�7!G,\�o"'3��놝�)5H2e2��a���9u4�3��!5 8�xVxq/��˼;��G��`�>\d���
�W����FA"{�f�jO��k45�hxh��>u�P��������G�Y�L�����APo0Z��9c���(/�e�갲R�h���9�&S�>���;�G�)�DBP�=p�	^���:�̤�}�M#A��z��.3β�j{�g���@}�x�xԩ9���I��a��=���l�H*��%: Z�>��o;]s�5��2(��� B�����3��DT8�44���^,V©N��"���y�Z�>
�gv�;���������I�#��R��''�a�2��k#�i����'=�������
��蘌^T&�H��*/=�N��n�R��SO͙�	��J��\���.��q=;�#����jw�N���-�>RhIN�uVݷ� AxpT
�1ֆ��p����k��f�ޣu@i���Z�:.ue�.��Da��brωr��Q��q��q��u1­�b�AX-���]���h�/�}��
^��"(:+��	�Ԗ������@��B����#N��lZ���S�X'�����@�5V�Z��г��5�yM^<"	S�i��#yP���0K��4��[���wY��XZ��KRJ$�v���C�$�[B������n�|����f�\��g�s�q�\Cs�[jw�"4����?�fAt���gW<iߘvqϬE&��<��('��Â4���"B�Y��#o�02Ȕ|.='�(��]5�I��J��n�E+Р�˿� �IK	E����!E���s]ų\�&�}Gu��q��|W�6��a���;��&�Wgk���=��C��S�B2����燫�U��+���t���SdZV`�l�O�}���$E;߯�SA�A!�gGi���f^��G�AEY]B�8���w�Z����6���;V���@����pҧ��ȭE=Iۍ��;d�1���	\�E
o������.��]_��ɾT���᯻x^��ԽO��@�1��<�n�����xĥ�D��k�ߴ6+���,���@�a�8��7�4Qf[��|~x�J�2���e �4�g��ѩ�]g[Z����K܅��C�A��W���'[�� \e��@��G��r?Ti��~�D�;[�ǆ�|�̻��	�!�L��m<���P,�ǈt⺪u�_t�D|�d�>���[M���@g`;�/U�:���6�zs������z�r#K���cq(���`p5jG[�
HJTS����b�z�$%��-4��6t��J�������#�m���
������B��5�C!��A���2-D�V	��/��߯q�0Wo7*"����?r�oi|��x0l�����v+g����gd�0�E5.�(�U�Y��6A�z���卣��pBq�[�eF4Q�Kv[Un�D8�;T �����,�X Ti!�#HZ�&,�K�<�u0J"���K�� c�v�!����y��!E��W�m��|5mA�𝌸Z]}ʺ*1~b Q��	�Sv�]�F%�Ҩ4���/�q ��R�8
��Al�M�#�7a���0�Ã�ɑ�>�+~���~�0�����������9���i�<dF|�)c��R���f����s��q���G$־�ݙD%!I�l�or�&b��i-9��D��?�{����I8]�����h�&�H?������ 4c��~��j`壬����+Yݴ��z�lL	8|�SLT��}�'���H��������9|V����鳯L�! ��{��������Mϡ`
*�e��V$8�O7�=�g=3W;���Q�M���3��o�R�,�>p�;�xS*��g�^�j�g?���ѹϰ�0�ik���O��p����]��f�V�ǃU��'sD���{�=����Ue�±���-�2{�^H��� ۆo[���m�����+�_��EAA^�U
�����!(ĿBӯF@^��?*��紉�P��:)��/�� ~����n���N����öQ�*�H�_F��}��!,���bw��Wۖy��}deQ��\C�`h��(���+���_l�N8w�Sد��E�6��%�6�e�§#���_K��R�v�O|��Or�?���7�-�a�*�z<GĹ |�BL3��D���c[��0�u��#�������!2��J�G{\\\GYY�ί�.�
T>}�lE�F�Iʷ?�M�N�o������$���ةA��E�f;��L)Y�O�a9�6}w�,��on#�\�P���;P���x�����/�u;O��ZC}�&�~�������;ym=YHZU@
��y���NOG���2: ���̴}�v�6��7���"d�(#���h�&Z0)�X�_��v|؄�N���|q0�T�P���A'`��0z_Sɻ�X���C�f�m�����
Y븀<��̠n���t%�	���d�A���)/ e
�US��������nMYz��v���Zf�D���s �*p܆�n��]�N��p<��� �����]�Y16�OpQ���.OIl�sM����п=7R����g�iv.�o����}b�gr��M����>��C�i�mq��6�: "�ɢM�jVH��,�}&�f�H��	U���q�]-���͉��70s8�%�dq�+ű�j�XY�x/��5m��;�����8���������?��B�ѝأ�yI����"�m�y�r{G{�?A��N��}��^3eR��"q�(t���?hP�U��a�&Q#3Ħ���E�nN�x��'v�&U�۬#W�Ϧ�\o�sa(�k�Gh�O�T�QWS2�Eb�zB��c#��$C/����(�v=v=9���u�Z1���G�Znj�G\�Yp΁��wT��U�H���:�#�BP̟����C�D�����u�׿v9���F��G�U x���HV���j\WM��a�-��G�I��Ԙ��-m��/m���UP0v�,z��>a^��Ⱦ�z?ز��S��e��Ci�ĜK�4p%]�N!�d�Ϩ�BW ��k�����(_�V3G܄)��5�Yj���!�b|"ѳ#���UTTދ1��r��2��kP��N�i޾�$�I��^�A좰�.rf��`��8i�*!0�y�?X|q��6�IɲV3��{��O�������y���x�Y%���=����FoZd?K�~��
�����C�����{A~+���5ӂRw�ٸ*�F�o4�7'�{ �{�N���Y����O�4D�^��c�y���"�Ju9%W��ra)��]2���z�!��D��Я0���<�x-�ݷ
�3zܐ|����Wh�x��\����D���J��AyEx�1@�(�q�c�1�C�[!V OK �C���*����P��И���z�� >.�ht��R���%^�@ no >LE%��d��wx��<�)N�y�04>®�|q..E�I*6`�����(�Z��^k����w:�Yج�o���KF��-���GP�X�uM�c����39@b�����=��� ~M��G3�l�?�
JX����"��5��ʡ�w�vC�&!�2��Yu�����wһ���j�ޥMoy�/�� O*J��ts�x^���(l�������k���.��������Z�ގ���M�%4�3�p�+����c����}��8�����µ������l�q����Y#�z�X�������T6��1S�������g^�u��j״�a�_i2�5&Ry b8�?���i���QLݡqn	D�/mZ&�3eS�zJ������;7�<x�N4�Bj�b�w����|
`�Y򐆈~�!T{�i��{��]D��.ɼɹ�zZ+���!�"aJfQ�}��/Gc�lAP����Fc��%���y�ڀ�����ii��l�7���SE��;T��Z��N��p_ޟC����x�hg���J��m٥�;�qr�R��e-%���xO�Y17"h\�F&����:�.yT�?���Я-�K�S��'�7��
 PQ����#�Ty�9���5PJ(� �TF�����F{p���x���M�[D37~�i&��'��Mrnʫ�v��B��7I��c�ޒ���_����j��j��F����}1�`�x�'�v8W>��j���2F�?
����
FR���h;bo3ڀ ���wjh�m@�yS��qV�k�;��2�m��1���W1�p�����7�����8�K�۴���&�O6�/��h�f�����<����}Np��N�yh���9~7
y�nM��.��K4�Cc��_F��Å;���(*m�^|�}���2��;A>Ç�,�t�a�s�WD�EB<�� $�(��^c2lyD��5�U�5��fW y���"�quޯ�+s<���A/W��֝��3ٔ�5���p��Ev�ߌ�^�TD�-&=��+%"�k..�Q{/��B�� .	���"��˰�D�һ5�W�1��Bbn��u���{X���rD��o$�t64I
�pV
5��ж���Ñb�
�_��'}�vd_��2��|<S�Bg��>�HV#���4�v"s2�g}�xu���Q�,;+�<5X����ż-2�* �jܒ�Xy�zff�v�v.B�>��3Z�}o{���*��8�z���eі��ڙ՗[��8�h��	@�@� ЙI]]�!�����A�g޽�c��#����#����z���VBՒ��]h�n��//��	>7�+(w6���ƣACcu$'=j��V0����&��'Q��)��"��6��0XP����D{��ǤrQ���QX��n��g����e�{%`?<+E�	������ID.+D�,d���պ�TF�^L~�^~�A��^�#�^=ZV�	O��pS�=j�DF���-�1X�H�I����#�W��PS1�����z��.��a�a]u�h�@���;i�.P�<Rx�>c�<rr���19EGu�l��X:Q�d���� ��'�Z��t�g��'1��?.T<��X�V��T&&�2�t����?W��kȬ܈�K�n�S�;y��>N�%��R�N�[�eL&�|�H�O���{�t�D�h��H��wyZ�6���T�)l8e�ǭ�v�ʂA|�&���Do@0�juʠhI�y}fja� G��a_@��^��Q�����M����E&}R��T��7�,L�pS����l�c}r+u�r�{�{�]�5������(.�&�ޯ�	�M`<f����A���Z����~{c�������	"'ᬳ}���67���L��g��ɋ�ɩ���%��Q֝�&;/��eb�m͎���ެ�WZ�5��?�7���|y����HFF ���>�Nm7μ�a�`z|GB�J��v��7�$3-�i�����m�4!�2��\�O��x� Aq�J�m��$ͻ"��+��f|'�u�
�6QH#j�r�QM>jV�m� �<f�b�w~.e�ёލ �j��*�5-.g�1��ss\:�3�+O�|����!L��K?�m��
��毉��׮1�q4_/�1
	�&���yN�,�%C�F#/b��;�b�`��X����I���֣���0SK�b6�p��a��0�8�/����w~��wL�y��5�Rgo��^^�(ѹ���:��I�[@��Ո�a�[�I�ZӨ������j*�|/��x�\�+׺^O�雏'���dф��ao�^� ��T۽%��An�������oS]�el���}����~9�s�f����!�F5t|x�RI��L�F��O%c(`��A�O��|:\ɸH���7�&�X�z5�R�di�$��>�6j�������s��A�$ه�J�{������1�<�N���O��2�J��Z�6u��񱝟׉�OA9��Z�����|��lط3S�(��ӲK�NMem�ƅG ���=�jX|�URr�r8�"�&K��\oU���XU�O!���u��(~p�PH�|V���T�s�ƚ?>����A�)w#����nԭ5����LW���z0�0�"�8{X!~35�����~"%��ӕZbU��.��3���eKC�Ro��/s�i��zA��j�]?�Z�� %eX&�b�
�֗�����8�6l��J��� %��R31a��֞�N���IT`��]��Ĭ�H��W�j�2�V���n�h+�.���7)�ғ!�3���4AT����&.�7��9����~�װ�Y��ʢ���ќ�Ƥ�B�,ee��@lWHj��mE�	��G��3�.���\��EG�'�w�o9-�0��s��{Z[��C�jh�w���K����S�>��an���3��o�o� �fW�^�	��d�V����R���<��P�C'S�߇B�lBV�p�� �:֗���V%or���mݥ9�]�h�y��2�G]qndBs��L�FO�p�G"*���5ǝ����M-��W�|S������\�'�u�BQ���t��8���pu���˽&S����q&5�v�����Y�]�'��Є�w�ʒ��l�L�Ge�S�����m ���[$�K1��X�Vu�ϖ�Q2�R�g�F�ކC�ّ���_> x�Y�p��ͽO����ș_���fLUhfH;V#I��[1�(���IM��˽��B���*��C����߄z�� 4D�葳���q��]G����z�;�'���.ݼ���ⰰ�HT ,M���`����O�f�V�寍h�6^A����(���t+2h�b
�"����_�!�h�JYx��W�ϵNyo�C�nu��>B,ۤ6,~;t`?���]����M@M]P���"x��ۯʏ�� t���T�o�P���3�����掟��0�1���tK�[�۶�Yr��D�~-B�&�T�%�u�k����l���IO�VA��6T��:H��	�?l�$x+Ov���e�S����g.Mt�3��K`ͥ��J�/�4�N��}0�{S��n�/��YR����� ��^���@��7y'��Q�T!��o���HU���3}A��d���y��K&�l�/��s�������5w@�[i���~�A��� ��,�3݄���	�6�f�M��ק�X<��m���~�~��X0J�{3�D�|� t��H�������)e����P��H?��O�$���g�>��o�oa��s���I���h��#��|��v�)1�,������;c~�Yj��}b�N���vK3��0�O[?��l,�v�T�|�sy�x���G"7�5)X�O��jf*W�y���ﭫ�.������t�Aliҭ+�&j)��1NB��((��=q=��nR�ɦI���2�rȲ��j&����I߸2gc	���������H�y4bY9�����(��w�˾�t��j���;�k�`dx+���{M�JT�������Z�l�t���|��t��\��&��}�i,w3]�c+��?l%���m�b���9g?%Yv������LV�Z�HϬ�^	d��������j�J��k��x]�E�n�X�E&6c������DRZ�i�B��S5���ug��Z��'h�NN�0����4$����\.�{ށb�i���h��
�Y�2��Wr6뎥$��M�0�7"Z��Rs4� ��Z���O�88%�ʫ:�����4� �g�g#-��ڎrӳܾn�Bax�iȷ����`H���ϓ��b��׷�7�J"+/0�O���N���AQ5j-�ž4��y��xQ	���$)��.�?�b<�2$�>a[g�s�����_��:���zZ+�8��g~k+�X!�*�_;��\������	�B/ �&��ө"���ZۂGנk�0��ڦ�_�KSM�`�>�n\�A$�mH��.�ؗO�C#.�AQ��Y��ZX��ug�<[;�ʴ+�?�Ow�x�O��VaH��u���⽈8 [觙�&F\JO��-�I��TӔ�[���E*�z��C @�	3K�>
�g��;AA�����\/�eԶt���F ���PmO�;�?�e�9A���o�ݣ��'rw�(�bA�֨<���Ű��	T���Tշ�sv"�x�UE��t�=�f\?N���KJ`�2�,5?���9������e)�7���P]�z��S���TAe{���>�{[�NYi��^�;8��D&��!���K���X�p_)����^��U|B��P�8�4��HڄT$��^�)<a]!A�7�QC6�������M�f���t�O	ib<�����?�6U���KѸ�t�k���`�%1+E3�`+1��+�d��xu���}��j���$�L��
lwH��IH�������5�=aݻYH�W� U���;�ꆾ�PE>%�*�hV��"L��L�K�!���3�}�C_��7]P�L�E����D4<+�Q��0�^yX�Un/��e@y͟o�B��V@���k�6�t��c�4�S�_� �!���(V�<��Mhh<s�!�t����$��6�L�¬34��$���!�'P�D��nm�Y�|׎h>��9��ƣ�Q	���5l�^͝˝n����*���M��s�y�Ț�<��JA���zKP"M�Mm���z�7��8�tA),@'S%ѕ��,*f�����^�����Xz�2�P�DT����.7(����e!X��ā����h��&S�����@m��Ra`����G4��	X�����썶p��[��ZQ�0�^G�l�E�����Xi6���Ե��a�"A�t!?���y���C�M��T2�]�6��"z��9�	xA��F��lq �Xx��X��2l�c�Hkƣ����5��3���.�J4��u�Z�����i�����]���e�`�*���A)/�@B;���H��9���9�L+�o�T�����B�f�^~W�I��M2��CZ�L� �U��E���dqM�&4	Ln=W`̮>/[鿜��2uqHQX��=����'�3����#WV���p��Q.���0�c����f�L׆�)ɗ�qv�70-ND����?_���oc�������+�D�5��'����V/��=�ً8��xy�=	ĿY�4S��Iω�ױ[�?��BY7�-�~6��n�lyv�Bc�pȹ�S�W=����t2	����hQ�0�S0�[U$�\���V+����Ի1�`��/�,y�y��,�.}b�ߴ��6e�@����%ˌ\n���,�~��a9ޙ]Ow�!�l1jN'}F6%ڿ�6�M��/��XU����Q��ʸ��\�8r�z݆�?Ӓ��R��k��3R�h>��'�N'�~26P���d�5�t���nL�uj�$g�q����0����E��]LȰjF�X��_dB�����K�w0�Q�(���/�m��y�uQ��V���M��Ѡ`-�1̏��/:��"c1n!K8�I��*�	5U�����l�L��w��x�u�Ug��v���VZQ]\'DgK�]���$�T܏��Zfh��U·�L�E���\����M,-�HӡtǱ��2c3O>�*5}t�SL0��'<s�hB���>H����%ѷ(�H�V�7l}n��XE<����~mx�n!�&��Nc��7����s�b]#_��m`���J�����(�{K�����6p�F����zv�������a������t�l�9�ǍͤUԺB�d��U��G@�s�h�6�����4� y��H��6��Iȓ}��ލMN�95��Qұ,\�]���fY�yA�������zB�I�b&v]k�=5�[�#,�^�(=IjjSd6��:�b�^S�RR����D	�~|��l�* ��!pB��h��9��A�ԗ���E{S��E�Y.lZj�H��-o;�8J� )��gL��$�8���D� ���X��o�?�?�����XL9�����'���Ŷ�S�5i��Ki?�b�ZʑV�Ϣ|�t�4N�<��z�|G�����'ex]&�V��C��#�t���;W1�a��֎�ݝg�/6�[O���}/�_�<
.�1�җ���H)P����i��-��t��Uf���t���.��9t�J������`8)X�i��F�џ����Ki��{�P<��o��@E�' B�H�k�|�?Fp�B�a!���鏟�1ǆ�{O����\�~��K��=E��B�AǑ��]Æ�=u9K��Ǵ�x�3�?y�3(�4�,��B��!H����H�I1�I����r���L��ڙh@��9�	�g�A!:ӱ�]E���"�����)FeTdZ`����d���xR:�\��me2��g�h/���^%�A�Vpu�"o���䉈�][4����X�l��ѕ7��qG�T�zd�$��|4="�wR6K��T.�c���&;�Y��xb��&*����ĸ��1:g>_O��K����?pg������'��:���x	�{���z��Ͻ䃎J,��\Ř�ңp�UL(v���j���7���$;[�/w1/�A3�lQx��������`%�<�/ey��C��_�� ���]r{�!ou���bM�%�Fx+�+��8�K�3�ML��S������h���c��?Ѭ�:�[�7�s�P��Bw�a�I���g������>c籋(tl��W��x�5�^��M����r2�Wm/ @�EU�-1��܂�r�ՐM}�v}9l�iB�P�1_^�ȥ�j�Z��+8�5�kW�5f���!����l�վ�ǃwZwY�eB���GH�%���A�#�<X�s~Os�s�E�Hf�!cL����l_8���
���ƒ.T�p̶����͹��UN�}�gߚy�&���%�F����Ұ^�Q@7̸�����u�X�Y����Ũ�y�T_�(R�TD���)u��t�!���	v�9��HZ\e����c[��>����uq��|(��iO!�R���8%�	[^���C�B&H��H/T��&[�/��Gmk�s��w}�N:�c����� �fIrZ͟�X��S�˫x��Fep��'�� ��r$�#��H���Lt�MI����r�ػ�l	���bl昳\�y�.��s��%��a�젾!�s^/�J�V�ݜoZ'
�;o�{��a�!(�MN��I�;J�u�X*$S��#�/BF-��t���˂��cg̽4�y�d����9F��2[_�N�j����c�ź��' �k�EN+:���v b΃��ƞ��,��C��䧺���bR)����]:��DV�2��<j�3+�}��V�/���.�)NpW�����y��G�|��kևю^���jj����"���!y��h&N�T�A��aL����Д��E�M��k�Q�	�ma���ȷ<Hm7ٛ��Oܨ�R��w`��D�yF��מU��X�2ig,5B���Rۓ:e���3p�װ�y	�TFC�otJ���D(Cu������`��6Ԩ6��w~Ϧ���\W{�IT�|�5$\�֜�x����%�l����3n�9]�B�/�[�au�����G��W28ԝ:P��􀲿��dv=	(Q]ˆ�̥�|;#ЛG�t-hw����"�,��ؗ���Y�!��(�+�Y�O/T��Td�c�����V|M�*^�Z�OcJSNo~i�'>��;T��;�ؿ<BF��j�@��.�1,�������l۫��2��w)k�jٿ����Mg�7VOX�)_R�p�<q*��۽��K�������:v�댍>�%)s{��8R����א�
��R㫕�Ɲ,��.��!��t$yfI��y�)�ϧd����H5� y�/��"pN2�z�jF�D�^,���;�G��#�|Z/��q�Y���U����8"���ЩA_E�Vʄ0I��ʡ��V!����c�h^��������9"�1�NS���Rʤ�Fqُ�� �����b'[T�W�)��ʢ_� Ӏ#)щ<�:G7 '|�����&�T)�G(c��nZ|�����w���g�o��T�6�~X##�3�A"�ԣ����%�W4�/���E4Zwa3*�� �T$I@)}s?��_��h�/y�(HߍOq���6V4����r}`m)v���$�j����f,�z��؟�ǲ�XYm�y�est�oLdq��%����x�˿!�Ϗ�h��E��ͣ�B11�&Fء�i��O�%��]����R3�
	�<T{�k���ȭ)Y���%�l!]�-|W�"p�{�AL,~��_�s�\~4���e����{��m��-#v�!����Y�!��{�(��|��&�� W�U�I�nZ�� ����;�������~#i�Mϵi��bfl�-o�>K?)���$�n+��䅴������X	��L���A���nޙ��Ɓ�i��N�X�mk�X<���+��v�;b���4����S��>�����=0��I��@H?K�D��#,,���T�TSe��m�[e:`HX9��E�<�K�@ĭ⅋O�[�FJF�Yp_!I���E���i}d
���qd ��MSD4c��<	eT\*�
<��qC(�I�6��(�R8Ii<�S���w�|8Hi}
sA�CF�|ü��j����_��ܣ��A,��]�O��*gJ_������b@N�5��1d�e�+���M����1/!��f���O8h�)�G�N�n4Θ��.^�tVԬ��C�p�~�>�b��ewK��mL^��Eﳆ�~̺W7��o��j�?� o�F�q�^Q�P)G�=��X.��<� ^C94�5:)�*g�s ������ Kx�X�e0��XH��!e�j4�߶퀐�����Z�ttt]3JfSi�+���V/?��tq���	[&��.6��:��_��o'��->�3	E����N�e�ϫ�S;O��ܕ�ʰ�K�|5�b���P3��rGB_���W�&���o�r$�\!��]���kF�&&�%�'2`��5j�4���E���à���K/di3-N!�'�i�nRaf�;��/���;p��}�����^SU.�6���:v"�p-p��%�I�x\g��Q���G-�eb.�M�Y�'q,���wj�Nb�9il���W����8�1�G�V��].�_��mSs���h~$��+����BS� ����٣���u��uY����@ $j�N����R� �c�\�ϙA3r�/Bv���(��p�d.~���l�Hd���*�?��l<\���?��:4�k��'�[�t
N�����!k�9�`��Bԋ�E�NZS��Z��
�Q��0ey��]�n�UQC]I��~�Y�:���Z�e+���G�z{��BA���x�%a-�����7�,�-{�����>�Sс����@.OQ���"�ߪ��GL�V��Q.X�6,H�E1:�,��?�]��n̔�R�SP �H%vˆ6��eF^����=��W�m��*{#�I�Xb��>�|ĭ����wa����ED�ȫu[\����*G�Gv%*mkΕ���O��z[9���h���tFHy]U�=#ַ�Zg���mVW2�A��Bر4�)��W�tUH =�:vGySd�d�8*� �bb;��;��]���!�6þN�m�D��U���T>�ƃu�	魖�.H)nF��)_�x6���3�
�ztu��vq�(�΅�Y��^Uf�g���o��L����5�����
�{6Y@0��WKc'�sE{�%�s�������� :d�]���P[ύ��\�R�M��-�Y�2	y�/u���D�Q�hW������_�J���bF{�]���>'\��5`���&9)Z�f:�?a����������5C��D��A`2��&������R+qki���/j	�b-��/R�\1�O��m1:����'\YH�>ݑH���͸x�K%��ȴN���pI�khW�Ib�O��"̺�E�_��kG�k�%�����Ô��b�Cz���1J�:z��3N�h��w�{��N.�̮��>%6���(�k��p�HK����ƜgR��gZ�x�)����(�fy��/������T,���e�Nm�|p�v��9Gz���DW;�T΃.R��	feNp�2��N�Mt��\�"���[�����X�"M���Z�BZD�pe�sm �"}�j]6���|�IJ8�:/��t2�ϝ@Ԁ���6�p��@��G[@x�b��FEO�����lo��ϒ(���ۖ�ޡ��զ�ºoNcޓSS���WW����wȧ���Q�F�����⨲���7�����̽꽗E|�bbyxsH��wZ��J���̐�(�O�ͼ����`��]�en#f'J[.v�l���XZ�4:u{Td�8%����ɪ-�-~������]�dLo���2�D���/�B�����E_c4n}b_�=�����,��mw�!�����D=Tob��kj�-�|�>�>j�c��M�d���^r7��b<K<�$���N�p>��3�|�6#� b՜��yጘ��oj��pu���'�DmP�)�<�|i_V<K� C��M�����-F75��3[AC7�%����L=��p��1~��s.4�۴��2��~�'�Jw�$���S��.��E���W�NJE�1L�=��l�x('j�FD�w2d�����`�]\�9��bAg�*z{.���JA�Y�%v�mk��-�w��J�ۚ4Ka�
��y�7���z��[��R_$�s�T]�.1�{��kKZ���{cq�r<�KC���(�.����A�F�`ơ`Q`�7�A�z�+g����H}Q�G��* t����6�R1��(8�~d��������@�@�$���B��q?��7Ñ+{#}�s��+� ��И/�7���������/8q��=Ƃp��u|�.�i����.���#��Z�f�9�@E>ȗ9Z��;W��	
�&Qx]@��΄���<�]�!��,X+{҃(eS+�l~?�y�1�rGEW݆^�??�@cLLP�0$"ҷ�?nrDML��H��e.�A���W!�%�	k������Oc	�x�B�u6���3��k��f�m~�[��'�9�",�x,�����v�q�.-��g�_�c��~��k�"��g�l�}�a����Nqh�x�g4Й@����v+�p���q2VJ����y�<�~�3��ѫ�pM+w�p�B��_^��Ā)WK����MI��I�>�"��⅛���׵$P�>�4*Bc���nL�̎�t�F3�6*@(��C���� ���䍞�|��7Ѳ�1ZԂ�[�_�B8�I%j��*�&���P?YT\��e�L�u�Ϫ��7+P|"�Y���W�v���zx+]�W)�h[�1��ܕ"�����(=��L%����y�ɀA]�OM8�	%q��b2�i)��
����8R���m�V�@=��z�:b��=�s����@lY�
�TR��<�K�`�����`�h6�]�	|Y��|�0�?�V��!
��$n��n{��P���4�㌐X4��R�o�*}WLT�>[�����ۤ����%5 �21�v7�;Y�k�f��@`�J�9�d�Ǆ.��|x����s�7�Z	J�t=fV��5b�;��(Fn��v�;g�@��0qݤ��Bd��;�M����|�c�O��֑� U�@�\,V�d��������A6�z��Q|�ڪN�(9�f�Im�Nk�j7�X�g��M����B�
��ڠ�"�7b��:��J�AB�{�=���ǉ�ݵq����c�$V/��J�pŇL�琖o���$C��s.
�ۨҩo6@�4����sY�Y�2�笭������.w�)��ꍦ@Jl�ݮT�M���ݣ�n��	b�p����t�nt���>��R���.n�U�� �l7�A��a�`I>Č�˻Cέ�2�n@�o�H
���|��Lk)�8Κ��"��}Mڬٵy�1�~�S7��{���\���w��������,4NM�_qm��^>_�U�Z�Y�X��l��~�d��tL_�iUW��w��U`9F�6�����qݨ�BaG��ғ��d�u�3�C����P�6��J�k j����ȓ�kg�����8,�Rx;� BG�������R���B�hm�nE| /���.��SSSN=$��_�b߹w�
~Y)�M�B�κ��ܨ��?/�O�S�s�oZ��AO���W�^#ܒU��3��:������G�fUQ�M\��,I�������-y���%���?�N-Tnj��7+7�T�7�\�v"d�ʊ
1f��v��uS,f��2�o�.;��͠`0L]2���+3����.�B����L��J>i,�U�����/dKA-�v�����B�I��
�1<�^S~��N��=�/à�#��N����O�\����Ь ��xb�܂�٥xP�{V������I��������SZI�g+n��1϶
kҠ�)q֙�]�p4��-Wf�o}ī!��WEs��֌sLE���L���2A�FD�ٿQ�O45���^�Q�L��i9� \Baޤ8uW��L�s�d��qNUS6�JiTgT�ܓ"sa-XTOˠj�L�@l1�VH��	)�W�ΦD۔�/�lu�U���i��"4���SB2})`y�Hl���Bc^V�<�cpJݩ�`���}� c��c˚��7�S�BI��"NU�G�\�VQ�E+��C��D�e%�qz	�^;[v�3��I�L�C�q�YHf��rQj�`���z?,���T$&�M^{���n����s���E���B�]e]��/��}i��\��[\����*kE���B�mcG>��D\.s�H�����P����u��q�mAܵ���)q����-պ�M�����q���TP�;���ʝ�;~���)1��)�%������3o�֐m��}����#wO�L��� �vT�~���		��? ���l'7�W��2 9f� �4[b�z���)%ԣ�{I)����� �@]��#������!�-���J��c�+�%:�m��f�(ez�ߜc�YвV+>���s�u�fn������I���Ul�P�)�ǋW��賰_�2L)ʵ��Q6�Ax���gw�	/���M���C�ݓz�L�S�'�x\r����×f�9�a �Q������FC"A�N�b{�=��M��`�_*�eD�[J�S��Ԁ�Vdg��9) �EG�C�ފ	w��eAF�a�I��!��� k��35c������D�k8՗	R��;�.��b�ڊ+rrl�Р�
	8?��g����x�@�)Bl�S�N8!�?Lѕ�0C�Ĺ>�KN<����x| �� �+^������g���6�M�Y��0Q�����we�Z�@�0�
�yӛޔ�w���纍���u��s�'�9�~���W�����`�����1xŊ<��L��9�Z�^~�Eu���r��}��Ҽ]O�/���ݕz�V�wݞC����Q�kH�@먭�FO+�� �#������/~q�n��D��Q�
XVҳo�]��Z]�r�E= zjq��1��@N+c�� `F�S�=u���q9��Zt�����O�Ld*uۉs%^�v��d���Tb�Mh�Ü�!q��Q ��m�C��0$Y�\88����~zf�_|q>�{�J����ʤ�Y& C?D&|��_����Ȁ� �q��B��b� k�<Ϣ�Qv: �C����_�>K�<����`�1�'�@�K�ӷD]�<�(�L�����!v�$ �Fθ%R��aׁ0Lx����h��=5�gR�#*=ݩ�ڗ�w[c�*��2r1mrT� ܞ�KePpב�ȱ��S#6#��T�
fZO�0�3U��t�i*���L	�Q*�ؐ�T��
�#3U�3�2��Vj�v�H;Lq��Id7|����wU��{�Ȅ�n�^�|�3�fˆ�@��9�����$�=Lլ�� ��3����͟�ɟd��������h7���p�'?��p L������
�I��rl���r��Z~ٯDCv\�HƫK�2+�`�H��"F�dR4���Mg��9ޕq|���s�,77���'<;�Bݩ��|ڴZ�.�#��~��[7ϫ��ݖ��&s[ޏ�]�)I�49NOdU�21�����kF[��h�TH%`d :�"L�LQ��Y�:���0�9��t<^GpSs�7�8E��c]�n�Yb�f�L�>��U9Ǻ�םj�Z�2�O��3�,��M ��h!.���`��:�b�s��p�3����&�L�Q�����.���Mٜ�s> eyZ�O$��K� E�J6:�@���;R�%��Y�83^)��Z:�xvC������F����\���rD; �9G6ie�����t�v�:0S%�6�{��QV���e���eW�C{b���vU���d:Ʈ.S��og:��:y\��V��} 2��ѣde�X�W�.d��	q;˽L��i��_@f��l<�3��,��9ޫl��g����8������Єa�0�hw6gu���~�j�e��z���-�	�@�=���.�&6�@]M�c��ϻ�p�C��e����jh�:�D��||+�����j�[��s��Ϧ�(�	�o���|*m�
ǲ4�5<���'\�����#9R*3ǃ�d�ѡ�wesmw}q�pDs�����ɮ��+����eH"�>��@x�W�Y�欎�������m7]�J�`ٲ�/?p4��4V�9 ���ifG�*owꠑ��iL+�a<m�	��ɴ��9����R�w�39��X���Fd����9��3�@����+��e�Ɠ�{v�Fv����b-����J���m��I9n,���~�}Fg,W�]����I�^$�)^�N/PD�HA�qz'���1����=��bW�^f��ٛiVciP�-_��h���>���y噒}(Cd��i[ATPҾs�/�jH��r�w�R�Rc9d����}#�R&%>�,6J;��V��?��q��LR��Y����O�]���p�#�n�|�p^���1'Ǉ��3�&G��:T՝V��S�q	�g����f�i�H�S��2�3�g��_�~��h�ZM�:y�v�S>��?���.�I�2�`�{3p�vY�q���t^�R��ؗ���<I��x	 �|Wէl<�|,K`��͑��s���f�`�mF0zw�R�̺u�N?��#o�H}��ʲF�	�� �մ��E��)�^RW���E��hd��v��Y�x�*�����r�:�SnU�~ou�V�G0j����X���#j�婴���-@Ff��;2j���Z�M��yO��+���X�0������3<�(�,ʤ�2�7��U�� (�-�c��s��n�|�p��ㅨ��2>��SfZ��y+�G�h�܋�1LE)BQ>j]�u�V�G���j��"�+�ɛx�`��f�
|Zw�f�<������FS����Rw*l��L���7��T�]�����D@x�:δ���f�QS��E�7c��]��}z���-���c�N�X����""A���N�v`�ʲ�x���׬YsZG��	/������/oo��;;��c��Z��<FR��]5`����`#����>d&��d!w���ޛ�Kz�����=�<d&$@�à>8]8W88!��H!�	(I��4�� �E�0	����9W�<xQ<�	��t����I{���ߪ��~�vU��ݝ&���~�v�7�o�w�����w����C������Nސ�{��4�?���u��Vq2Ĕ�|6i�B@��^����`x�&.;��>y/jy>c|v�t8�s�i�u�F(�Lޙ�Z-�z��R��J�Z�>z9���8.u��aWX��b��vw�*��6\)�B��w4h����� ����;A��ױ�;󌶣��+l?PF��ڽ�a[)+,�x��ږ7��E[�X��$>�P�U��;N���p0�r8�AaP�;��fo�?�~%��ˤG��L��a�e��!�JNpƮ�jc��_q�[�V�;kl��OW4f�&wD�I�v��A��{��M#�+<�Dt����r�2��xm��GOS�WG��6e1�[�v���	n�;��C����QX�������̵��8ײ���SO�N;�����9�t�DHT#��6��T��z����2�;�t�q�{sv7IPt�YZ��M؝��
2�����בN���j�2��x~l_;{���t�lo��{rڹ׋$"��*��vsH�bt���k��*�����Η, ��6]�f��ދ���G�T�h�����L�jc�����O���\����0{̭���?]�i��ARw��lg�n�j��޿�`��X5gn1CЬT��Y�u1�/�h�Le��.��iԢ"�Q>¸K+լJ����^�J+ѐ��k���wΑ��y� [��,��St)�n&�<qW�����ò�Z�m�W���w��q��2��`�إV3�F��|��<��z���w��P�o׎V;�z�Z���c���!��\/���{Q>�8�]��22m)��=��k,�m�Q)��k^[6(��l��`�,��F#񐱎���^�l�2�Qqb>�a���MY�{�s*�r�HHr�V��r�V�]w�UW�jI�����;n�̺R���Ä+�RzԣN�L���l��/N�H�#h��ei�y!8V���e�s��;BEG�!�d�ܨх�]D���&�.2i��\)�1�G�^�@X#��x}^܁,v>�5���#덁�����An�K��ۭ�y!�]/v�R�ee8?��^b;R'�(Ld��@��<Z,�'QI���c��K��!���ǳ �<ܯA OY��m㦗`��b<��B��s�$>�ed���G�х��R/r�~�oJB��ȑ)K�|^��B@z�AY�s��&c7��"P���|�dL�RO���Au�wl;S,�f�v��M���tZ�Z����v�EK�O|�N*m����q���\5=�'-_�2��-K�{�/��ǬLS�>���rG�0��Ep�x*������������.�hV&�����'S�Qʘ�a!4j�S��m�N��`#;���\��+�� l|�7x�r���y8G�F!����������EcLf�r��B d��c,ovfoԜ�VK�@-���mJ�F�tZ�Vj�j���p)M�v�n�<Q��R��g��ZKs�-&�Ʋ��q��Z8�>�ff�a�A�}�iD�����Bo�kE��s��%
Μ���
��[�Bd��3�+�[��a�ڼ�5�=)r�������zQ^��Pzp�n�Ȁ��00�%c�a7q��wq��{S�uAuKH�	q�l��v�Z�^��˖���8���K��u�KW������M˦V�5����^v^Zw���h�S�Ioy�1��L����l��	����IK47��7�^a� �ph��Բ��z��YfJ���Iৡ�%�G`���q�?��@б�.��>sv$��q� &�|@'Sj�H�����{$\���`��9���2�����K=��d�m���s�Lw�;��� ��	˝Tj�ScvO�4gR�4�j�N�R
L�?��� �K�T�J��e��)�jm�9m���|���Ԛ=�;�8;��@؝ǩG���DFL�b#�=�.��Z8�>�od@Sk�ހ�KP���~a�7����=�D� �;!G�9'�+j�(qu�m�p���ƿ��N23�گ�Z|�%���ʖ�CdO#�}�g��.qv;4�&�-�)i���C�R/�P���duR(�,�[R���sL��ˎ�o��S�{V��I�Ӻek��g�����J�l�9�l��
uD�*�
#����/�A��R1��#}�@�zq*�J�0HbM�9ݱ���0�0�s](#�I!H�����8g�w �IƉ:F��4�ܫ40�IM��Y2���:-�b��#��?FFbor7ctb��Ip���:w ѭ��)�k_��\>@��_�j.����G?C���g���x�X{ww��>�y�/��?.�����4���T�{_�vfS���Cw�T�ו��y�;�SO�e+Ҋuǥ�D-�|`w��W����1u=將����B;#O0���P�7o�^ �F]GF��ɹ��ljp�%���A�w !�ƽ��9�k�17d�K��#�a����e�l���	�-����}�k�@�?�����v��v�n:� y�k�naͤ�$g��@���7�Ŀ��/���u�s6Q8��s���ɓz����IEo��@��D��z{^d�⊍K�;�W]s\���t�=w�]۽s�Բ�43=��_{lz�K_�V�_���_�����D`o��N���@T���i���A�L�l�� [#_(�4�����Ї>��R�1cr�4�>�bg�,��Ʀ�0�j�AS��h?��?�wQ?$����<�0eư1@� &�8�@y ;�b||ϳ��]�ʝ1�5��n�������
x�	s`0�3���9i��N>�Բ�bq���-w(�g���Z�6U:�Ԝە��ܞ�voK��L�4S��wC�dT�Bڪ�Ruٚ����R�0��d�g����O~*�y`W�*2�4Y��obx��{k��`C�Y�\u�U���漋/���+z��&��n5m�?ڿǩ�9~W��N�y��6b ���������}�O�ց^!yzق�~*a�8��>�M��A�z����&������ۋ.�(��+��r>G��ӟ�}0��乭�a�T$_`�7���_n�Z�J�z���.wē6}��t�Mo^��g�n��2�RJ��~��t��ek'�?��?�;��Uw7j���ac&>ӹeY���\v� �mDu%�*�
�qC�#{>9":s��rC��h������p�0W\qE�����2'TР.���h����y?L���2���svW�%�<���tf�x���)����n�|��~���;5�~9p.4P��戈Nw���=3�3�} �ukW�jj�NcWz`�m����4Q��r{&����F�of~�rjWji�]MS�O�ם�Z��4ۮ�=Ӎt��@15�-1?�K��s�zPF�3	�ِ�v�=ٰ�}9��/�D�p�����'�5��0a�Jr��y�X����c�3F!p,&�7  �����D�6��3S.�4�ͩ��:����U^�n�����DٰU��5�\��i-���og��>���c�9����{�2�mL���� "ЋqǲpH#������2����\�iӦ��l�r�;�5۷���]_�K���w��?��w�ȳ�j#�QL���]-K��ŀ޳[* ��>8����7\$a��ѝT�<�Q�A��pܓ�`��@�k;� �E�t��(����.L�Q���t[-#�lE�ar��<��S~�2[�Ȅ�;����� � �lي4���W{�9g��kV�j��R}O�ǖ�س#MTfS��Y�n��@�E�Ze"��Ժ����N�ʊT��Ү���k?��y�� <37}X��y�`�.v�� a��QA����:�������b�N�	���{���\_�� ��7lؐI�2����� �eP@���r?���9���F-�S׀0�� I�B���b�S��(G?�����_y��z����#���1�K��u���;���hh��w�<�v��n�Q/������a I��z�D	ڕ#d�����O{��r�Q��S\��q ���(r�$�����1�"x9����սa�L��U]�a�}d�N6Poh�	:. Lgְ���k�M��e���.�4N�c� a��{Lx:��Yg>��{���r=U�3��Zy�-�$=f�e�<�f��ij�Ҳ�'�fuEy���    IDATjt���F�����;YK��Ls���ʏ��Ud�9����l)�0��Z���u��g��Äq�e�Ev���XU\G&s� �er�~�oܸ1�=y  �F��"���[^���~�ٸN�]���ס��s�6H�ֻ�޹�[����/2a۪�^O*�%c�yb���/]�}�KW���(G��Z�利5I&��G��x*]ȇ�� !t�8�{��g&,
tL��^���Jd�g� qɘ����?������KV��԰�);F9"2�x\����p ��f�6�=1^��	+G �c(�x�;�^O/�[��%�޶�0�VN�yu\^��`��3^�"���J��g���Ք��� �J�SOӭZ�\��4�^��Jiz�����S���v���j�?�m��� a�� �@8�罅N'�,�r0a^xA��7Оq��Q�X�r����BL8�����R�0����~{lSc�x���{�gF�H�����C�0���w���c�0��@��@x �B�:����K������ߗ��q!j��FG�h�DG4��R��b����3�<8��m�*��|����W������?��yGe��ʥ����p�x�2]EA�@@��	;"jx���"ƀ1@ga�(����a��Z9B&� g�#�ZV�a��.1&@8�NV�#�h�y�E�1=���rskV�j��R}Oڵ}Kj��@�5�Քʬ��p^�����J��=:5*+�\�H{�&|mᩱZJ�V�m�Lx���G;*���d���+�� ��V,[�`� ��0a����=�����*`L��Ӡ_�=��<[��1��g w�8�#���b	���w�0�G���g/{�U�~����9"t����w�ؖ[ߴn�֗���3��!G81�z��Q�T��dD��3q|<n�F�h;�c-ch	L�0�^A��R�V!��� LF��C�T�`b� ����
�v��d"�	kP��Y��݄	�LN��	+-��9�L��}r��4��)�w@���v=�K	
L�e�Tji�UK����?�µ�go�����/�tA���$���~X�/��E9"�	c�Q���)DQ��Z�N���	s���Q�9By��F�҄#����
��Ș`c>��h��-�&x�2?䜋a��r&}����Z�HȜq>K�;D���> �D�r�R�0P\)W>�q��Y2&�o�r��mY>��	+G�	�<����y�Atw�Q�o*
ed�a�0a�)uc~G��	#�S��-��&���l�P1hX/S;��&L��LX��r� ,�	�	�|E�ӯ�<� l]'�# ��R� ̵��N�9p�/f����l��gow��61��# �j���s��m����&<�A�&	O���=}�SKӭj�:�4��ѩQ]���X�=3�>�'�H�wޗ&�*Y
�kD�]�y8�� ��'抚0Lx!�s�	S�h�21�u��"fg����BrD$&��RL̙��? �L ���!!�� �=�	�Y&�g ��N���	D ۧ�=��Ȅa�BB��	wCtK)]�eo���x�8�kA
�_6]��v獗��~��k:��r�!j�	3� �0#��ZL� &���}o>o� ��R����f�a�R�Q�U2�Sa$�\ef��n4A���@g6�� �L�Ɖ��QR�����K�;1�=r�W���R��+>w��$%���e���_si_�/�gz&�zr�Yg�t�Ks�i�@��4^n�rk�|��	ۃ7Y� J�SK��JZ���4���ԮN�F��=����O\�vݿ3M�Є�~�8���]>+�	AXa��1���A�w���0�	h�Z�����W�l����8A/�&l�@(�/@� P�/�cC}�����%��`BX�K ��=��RF��sW�ƍxi��s�� a	~���.��%�n�d��7�}�D��Fs.k�G�X�k����w�9/֨כ$���>��E�;l���S:-yT8�'0�όV�D�<u����9Y�a@
��B Lc����]Ӹ����;\��o�9���c�+j�>����\ <#*�3�%��;�񎮜#t,+��,̆�}��O��O������"7�w�m}h��c��@0~<
���Q��� ��^���k�涛k�s�=���H�֯J�V+��{S��>�:�T���$=dI놪�"�Zf��jj��Ӳ��R�6����|`W�����������R�3.�E���6�J4�Ձ�� �ع瞛m���f}��`�=�~�d9̫@����*^��+%$J}q��r��r��/��x��!MG��^q�_��aꎸ}"���g��7�pU&�|@�Uϕlp���:+�5}vA}��_�܉I�&�ўMF_a�"��[��Vf�JLeT�奍��L��/a�s�  ��+קs�9{�����F��P4����T��K�g*�����6�����??�Ӏ�Z��!`иѭx�k�PG�<*�5T�����p���x��v��m�c��ѹ��+���3�����q�����3p�7#��z�wup�� v:	uI�v"�r�,�@�R�B6F@0�7��l厲wzw*wHu�L%�O�	JC���vzrn;uJ�t��.�)͗�?$�I�����gg�\�,'�!qζF����开ðW%7�L��Ja�Gam���{�mhk��[��`�\��z\�T�s�|��U��|����+Qh��Sڟsjȁs<��(a�+'�B���;/ u����_�k�\�?$��B&���	��sR2aޕ4)'�f����	� ����m��ǰ�{�	�G߻�es{s�	�	Q�'W��swo�'��< F�ȃ�E�Ӈ���z��X5B>�|�+�7C���Dy�T@9�YN�`�#�tw E����BY�{;���n���\~^4�c��5*#8�g��c�%ǚ��e�<��kG�<���,Nf������ێ欲J��;���r$L5�X�2Bml,��͜f2wn7G�3(3���R�CFo��vE�[#3[9uJݝ���rg�Tx^K��l6�� ����9��;_!�[��ڹgjF}�,g؏	��I�eb(	H��r�e���1#Iq�s햿%�c��R
�k�>��@�}�Q��s,�IP���2ǵMٵ�9��dE�"y�
���s� �sAl�ޭ�'l�믧�a���.�b�'\��u�-7_�n��,�OS��e*9���5��;�� L��
$8ډ�ج�4L-�M������H�{�~��,��Ÿ�[2p�<�09�k��w��ϡF仃�#�����������Ռ�P4b�se@�!2x�`Y)�@�=ޭ;����*j}�2c�Q����dڳg:w�����]�_��J�(l�����xNi鋏� 2���r7��lf<�̴�e��i�T��;k�ژ:q�|�w޵m����i[��AS�4�^+�B��-pm�%@�o%��mS����$]}'�<���8a>,�K�����9DGy c0c�/����"������[W^.��PO��sb��˲�񪫮���SNY���·�t��w���>}4 ܨ�Ҫ��U�ze�#����Dt ����o�v�cX�#G@�u�u�96f���e��m�y���hn��Q@ΑLY��y���)�=���4���"��Y3�]�0��s�G��2;hɠbB"�*0+KP&Yב	��b�֭�
p��1��m�x�,GĐ�ٺl�,h������>l�=�z�}25�����fNٓY��a�|􈔥�;�M�eE�q��H$M=M�\���i/�BU��{��s�;��2_�U�e��-Cq@�?���j>�y�s�9'�>Z,Rk� n����\�} ��O��&L}�f����,��d���F�	��c{u��+����3�8c�bLr������fn6�9N��/H��N���{`>D�Q0����o�[��u���+�뢱2�����?�gBۘ���'?9?)%��9%��&	���$`iL\�g�E���02Y��׭�ÌP�Qɂ��80(?Ȗ�`�r>��f"�y�^2�AL*{�;�ZwϹf���c��ɚ-�h���p� A&��[���;ώϦ�e,ԩw�F3U�D�/�AD�0�M5��Ko� -KS?��M��ڢ����� !����%l��%)1.��t۲ľ�v'�U��k��/���,- E�s=�(̗�)&�ɦ��+�����,�L�9��6�tؗ$�(��L�{�b�6�1�ܰa����~�]��<�>��n��<@xl�����E9�<�����֣̄͢��i�bG��#3f�W��ys`\(��a� /�1Ǣ;�-S�0a C��VrԈ���s-�@wD�����Fg��*���!���6��;��\��VR(x���a��L����>+�*���@�� �����x^|��k���|4��֟ݎ��N��8���gV��:�%2�l���}麉���C�8�AX�l��HF���CQB�]e�\_�I[��;��l#�g4�'��{�����ne�[��]I\��,_L�ﵰ}u�P�c| &���|en��}�c h��|�#�޽��� w�'�-��IY�񊃟�籜��Ah�!��,j`���6m�t�i��v�};��B˄�m�㼩ٽG��*�	31��lot���y�幹�A�҅���ő#dt�?��2aN cbε߄��b�fA��1�&�*�@�gu�ڭap2z��	|�}d��!:�g�3�\�<JCq-�����!"���xΑ�����!$�l�=J9�݂z�ϝ'�z�1 �;�ZBjH=�!�,���Y~�)�~�VsS�a�u�N��+��h��}ɬd�F���H��.��&���Q��DgP��^Ji��z�����w�C��r`'j���g��{>��ًz���JH�>��d��k0Q�¨�<�9��!I�I��)r�zDB �Ω���[Ǒ�Y/Vγ�l��ԽK z}������Y�����^��_OG=j]�7�R9O�,�D��+��y����	��0q'��s����x�.�O�8�1�]�����OF�ae��N����j]�!�ݒ����Ч���9�#��=�%�3�D�����' J�	|�A��'+f���$	��`@l19�9�9���A�_mI,9��7H�׿���9�����7.=fb9��LL�q�?�*S���Lx��`�x�1b��{dc���Y9�	��^3�?�����+0tm�;�Ły�\��
��`���l�N����?�:���8�4��Xc"��D��`�C��8̤��_�vԉq�s>E�2HT��IO.��M�6]��r��w�ly}�(V5�	���W��g�˫�ƪ�AX�(6Ha'�tK��t�8b�����o��[���ԣ���[����} �V"�l�8���t������9�> ��~�<�w8���m8������E���?��qz�1p�	J�?"&8�����b=쨕+'z�b���w5��u���Qwo{٪��Q$[�	��hPմs��4>9�(&ܯAc��j�`�:	e$��ް�aF+yn���5�����}�0.����}�5Qx�R���y��r�����#��?N��	n�6�M��~���\'���W�XLTw1�I�-�V�W*���#�m7�q��-/[��G��g"��j���6wg>��n�[���̣>�䟫���1��� Ց|�{�a�H��s��j����`<�����|�����]]w�u�j`��������Z���A��z� ,�ᤠ��N"F�̶U���,q����	L~�zr�W6n���%�# ᱻn|��{�z9 L�V�� a��L{oγ2,Ns�0o���9���+��V�P7f�~?21w ��=7�n��*�v�;��v�wys���q�r������a��;�j�+#�\�m$��(��|̓B�x������L���x���	��[��֗?�)O!��ȯ��,���nٚN�hw��Y.�(�u3`��[�,�s<�ai>Le�����1C�z��O�3�ar�~����(�@W&�pO���y�AL���_Gd�Ca(��X������g���ԐP%�w����3���?��������֋9�@��SO�:�^��A���ׯ�~��W6�fb�ݖ����Sg��[�D'�%,6�ofTn�+��=��w���T������[̳<���P��@\�{~̝�x���=����l���{��#g>���R�[c��,=Vف>�*��t{@9���k�S�ʠ�)�r��7o���SN9��Ŵ�� l��r�ZjV��)�R݅X��������X���`�����KZMFjK(���[��:���P9b1��	ˈ��b�q��A���\l{ŕ'��+5e���D�$�i�{e��_tԁ�ㇳ5��`��A�\��W]u�yK�y�ܭ7�~��0��c� �q9ڒ��\��s�6� P+��$��A&2�f�{8�ȽnE � �� .�D�E���8Y�jN@��f��u�����)��7z�#	��M�9��;�a�Z���j�Ì��uy��/���F{;��v�#W?R�k@Y��t��#K!y�@Ў��
eCsK�7y]ȯ�>+�Ҍ�in�w��E�nQ4*W� �,q$c���0&���,.۞�(��>�F;r�!�m\F���6B�g$i(Iؗ`����0�o������谍>�p��(���9���(�H]=L��+f�1<�p�d(��G�ɑXd�Er/��! ,�XH��VJF&`��y!σL8I ~�0s�-Yt�#Ev��8�r��0� L���y����g�0,@�\d8r��8�5Pd��0L��~��v�1�v�>$�1��c�̎7l��VaE���U#$GT*��]y�/;�.VZ�ճř�@�`�	;��	�9+G�	��Ȥ���!�mGnv��� v��y�a�h����!Z�u�
�醝.�$� \.��f���K'��	o}q�?���F.�/c �����_�żݒ��ѥ��@8.m�G@xXm��P�@�s���� �0a��[��;�dA�/���~�����!?��s!D��k��D$���	Ah��u2�c�ڞ-�ɺ��6&H���5��r-�0'�L>�;������ƖE�^
͌k��刻����hd�<�Y����[���y7�
[���.�L`�bbr:>�Ƚ�ޛ�u��s}��VH���7�t��`�����{mٲ%��|��e[,⹑����q9�^�B�R�~u�,Wsq^\��O/-ڰ+DM@C�L�+������ص[w�)�p�B�MxII{p��?�Wd��X��.}��gQ�I�e۴;OOH�LܐN�ܾ0lb����b�PW�@������'��S��T�KʱI�a�&'|����`"2CGgwדN:)�b�c���W i\�]��b�<��>��d�@��k�f��ʕu�����Ή���!7�i�������H?��?���_�%�n�S����1���V7vV�Ϡ�f����|�K_ʠ��I��^���];{�3��@�\}��Y]�'��C0����֑�� ����]��^�i�������`��D�;�=Ԍ�e�
<ĸ�2[���g�gyt�W~�~!GY�C4��5�{�����ڇ�T1H.��}�W.]�G�!��H؋���җ�4���+ۨX�	&�C�@0�������{���
�H^�WdVH0�w��]9��k���N.����Q��,u�cZ'q���԰��ߣ���i�π�Fa���.|Da�,z�=��[-]t�E�q�{\�A��g?���c����3��_�u����s];����w `�^�'���9>�{P=Yp��r�D�@�h���҃���U����3�*��    IDAT�SG�`��8�/x���J��|����y�>s�"~�gӞ�lL)�q�^{mցy.�����y��;+��>�����g�4�m��詍b��# ��L��Hq?1ȗ��e�	c��: )c �aN��3t�p�]�I'g��a\�}�{_ޠ�� ���
p�U���5_d'�Q��X�����2b:��Yf�Y뉎{��f��D�'�k�젋����~^��^l�~��s��l����[7$m
�������K��F�SIF��͠�WN�j� 4H
�*���U�
S��?�4ݿ��X����yW���-�{CD(�r �F��`�\�m�b���p ����R~Ҧ��Mw~�����������?l�#��&�@���8&�KÌ�&Ʀ~��adweS��i��?~�{ߛ�p��T+���<kT�AF�q��s���b���xc��S�_�T����Ox�2����:0&�*r Mg��;���5�I�y�c���|�A�B�zի2���������|%��;U3�������������ۜ�Q���m��sd�QۥLN��[���ҫp�,z9���l��MR�h������1�K�,~.GVjRb�l����� �̄'óAF�j$:T�;<�6X�s���W����W,Y*�G
cl�L춊����g�O̩
*���B.Ԑ�_�,2C#G������<�Ą@� c9�X��ʢ� LP�e��b�D���c���]6���>��Ol�
{O�e�����ԑ�鬀��/ǲ�9r������=���;rė���<ؙ��zg��nY��A��p�a�T�:�5~�9��b���.�E;�����W�-j�Q��3��('0/������� ����dFy��(q��w�v������o���F���Q����Q䚥�Q�5�K��W6o�|��S���!a 0�3�8#��I��[tCuU�����	�2h'D���p���ja\SƸ�b���9�=a�L���fi��놌�  �����0B��VO�s:$�#�L��(��ZL�!Gp�TF��L��q����7�1�9��������	�V��9ka�D��AH��`xb.���Aח�r6C�Q.��N�ˉ��ROFQl�Y�zV���v��6�F`�w$5'���<��z��ȤeД��2�G��2 ��W��%H���C���ny� &ܚ>*�SN���m���߶|_J��S���f�y�]u{����-:�����Ё1:.���ݗJ4��A� �@t��&�@e!@LGD{�����g�� a;���� ��_��E����#��֕n/�&���d�H	</� +tL)�����6˶�4�7�	�3�r���|�#�,_9F@�ikt�8�[���A�?���@�!��O��Osx���0&l=�~�!� ���w�3�atݵ�"ip��	�c�a< �w���k�ʹi��	��|>%�v!��y�(g|^�A�;v�P�n�t���Q��K���)���5�[~��uw�q����zXkֺ�����[��jz`)8����{;D�7�4���"�(�p7vh(�ݩ�;uA�c������9��>��W�V�	W4N h�����8"G�(���^���năB'�0l�PX�F�1�Q�_����!3e���o�g��2�
�<Ϫ���������8_�w�I��z-��;� ~��^7�o�+�№�ɵ,'�����p���?�=�FZ���N&qO��>\��MozӼ�<�~����0��'�����alOm�:����7d eҒ��|��w�ˋr	�9O���-]�G9�6R�,��^�[�@x�h��)�w&��pq0u��aus ���#��q��N?���s��<���5�0���� c�} ���+��vw�u��.�r�}[�w��9ǿ)|�����mGJ�ꕢ;�q�c-�Xi�� �����=��j[��O�
>$�����'Ot�aA�^zi>%^/>���x'a��a�D�7M�h�S_�E���l�)��wd�B�:���Y��:���y�[ޒc�9��,�S��L�B�����s$e������M���>��g�3E�0���z�	##`oN�E��{���afۺ�і� � l���7�Xwڅ �'��ڶ�@�����r�K6l��p�{��VP3���/@ ���Z� 
������eR^�cʽk�����0ꅻ��2acL
E��,�����)<��Q"S64M0��ו���F�TQ��������i�2>�z��B��MXu�yv4o@�mܓ�Q�P�����������/Lqnd�z%��Y���M������e�.��V�ݍ��H����as���� ?���̓�� C癉� zV����� �/|���$��~�_�'e��X�\��e�FNP��x�esPs.���Z{� �ddL�2X�p�R���.��g�qƶQ�b~pZ���7�{��;o�d�џ	G~�]u7��~S��v�0 �<ủu�
���S���;��;~�Cc 0����ig�`�w�V.g�3��Cc��I��θ�u	5Z�(�sm�=d�~��p�m�96���&<��3&���=�L�byY��=#X<qp����g?;����E&\�rw]ڊI?�vA\p�-b��vRʲ�@�2�6���^a�0er���9F�	����G>2ow��R^�-�ﬣX>b�#s�1�q��5»�6M��Q(�EmZ��kDy",�	�t� &���/��U����2[���Z��=����v76���Zٓ%`������J�c�k�ޣȾ�u�N9B}K@�5��0&�M&�p��H�x�f@6�������91��5�(7X�β���Ŏ;��
 Qޠ��� *���Y��9X������ d���� ��>�R��(j�N��J �����tz·5��Q���D��v2l�&����4��=�}r<���BR�;��@
�E[�ي \�+m�6d�!��'a���g2Yf�*F%$�E�*���]>A�ϯ��W�r�)�c3:�y�5�&o���AL��Z��
�$� ܝ�|�+�<R�I�n���N�Eᢻ!$���H:s���81' cp.���u�00\%��_��_�bp�Ӊ0NB{X�E�b[dg�9�Y�As�E����ɒ�D����Ʊ#PF�Mt������B������H g�yf�>�Iy�s�o� A>@X W"Xhb.��I�a�`;�vއ�b�+�㱄�!GD-1u��X�GT���g�-���@m�m�M� �d��0�'�m%4A��9ʤm���o��v�hH�� ��D�8����H���t��������HbJ������]�� |��/Y�c��與��0�l�{��[W.�N���I\;�n�t�ob�{nT�=N���ӊѐ�y_�E?�\Ɋs��jT�\�E1��b���#�.X�����ר{~��pbN�j��a�]��D�b���=��
��6�hA8ztN&�.����y���vz�Z�' #�������b]3P,�JF�MqON@��cT��n��X�e `b��퇁���֊ \�,�w�S����@��)}d697`���zaĸ����q1n��1@�xk0�f�&e�]B]����!%�9Qk���H�r���͛7_tꩧ�X��f a�3k�����ﾜ���D����{g_�Cݳ�a��h���}:�����j��0&�TV'��*q�Y+�K��K�cdE=�:���lK0�1.������jpAR�s��Nx�%�<(b�덢SzO���
/�0,�C��xQ�Pg��4`���d)��k��_	��Y��z�����;@�v
+���+%Y*�Y14[!��� ��N��z(��я~t�	��j���I�0:�y�hJJq��0�@38Q��-���9�F;pMV$���DB[uP���,�%�L��Gς�2QI&�G�&������}ǅ+�{�2������y��4��[*wR�\�����I�V'�:�<�Vnw�q�$/�
��o&�*�@�\�{��{3{zI�&�D��d�2���'�.ty&���ҁY�u�)�dŽeb1!T���E�w�f�����	1x�i�e�:7�M��1�î��w�Ȳ�w��璙��YR�ַ�53,~0p��0a��v�#�EpU�pr���dH䃞�`�nɵ-�sB����wK��e�,�!Ә��� �P����l��	�"���a�{���/�\�R`�N@�� �0���^i��IV�Q�ʈ��<�fFك�x,��wu�hoJ�@XFo"F3��\2�'�]�s%�+����磤R��H�zR |��͛/>� ,3E�貔V�}�4��\�䀵
����I�v)e�&�H�q����ie���S���Z����P��*ai�(�`? D�Ȅ� l�f9)#?��w�x#t���5��X���k6(uS!g��$�J���X���~@c2t�g@��{B�`5�ıL�8b�j�Q��<h��6m���O���~��3�p�,���gC�ޑ{��@�7,�{�"Pdi�8�� ��g���F����8�F#����q�!�D�VV�#��aA��A�:�^��#|�E��BC�U6
%�%�� j=b�Lގ�fc��v�-��ǹ�؆��͹A7����=~	G��:� |���ޣ҄�j�0�vW�7�r%�sY95a�N�u��*��\��.�J�J	�픺l���J�fbq��u=v���iPf�k�u��s�9#t}�������P�<��2��������s�=FP�ɢ�s d�5���\���ʬ�	�� �`����������5�&y�8�Ir<	'�;N��=����H;7:��td<��;qT��Ǆ����e��´1e�A�|G2(��y�����[z�ߜ'���Ǆa�k�x�`D�(��ނ^	�h�
!��KY��r�D�$G�������A4z�=Iw��2^c�9`�|ꌗsD�� ��R�t�[��֋O;���E�}A����[9�m˥��c ��Ċf .������ۨTS�\jͤ��z���U�ͥ���j��R�6ݪ��ک�.��c�fsY��^S�7V�z}��j-�t�Sc)��J�TM�TB�贲�� > &L�ct���/كF?�yR�mW1a ��LP��bd�fň`j$����0��)���f�ê�P�� �b�ѠF?� <��t�g�m�E���a����ׅ��ѝ�Y�����,��5�r{?����[zP���_?�L���y'�9�Aa���rϵy������d�9�LX��!���_�F?��p�~؛Ǒ!�&���'�<ϼ�&H��p�$h3�.H9鷐&���N�T�ߍz�9��c�)��ฟvUl�C��o�d��;фd�M�z3W�X*�����J�Ԭ�{R�wn|�����MscS7�'&��T���6Y�ٮ�ʹS�\i�&J�63	�+�����ޣ�ssO*��=��nWm��U���j��J\�ԕ'F�$��\Q���?��Og��I�/��8AӑV���NZE:SV���w��Y �(p��>�:�VC�]B�Ыђ18����Q:���֋L�2z�/���(.�1M�ɐ"���m�l{�e�꿾`�C�*G ���w�Ű��ʄ�7��A��0<@�d&LPCꢎ����Ya�c�鉆pBU ���٣��,�~ �@v@�brv�&̱ڇz���ԍ���^��� ��7e�c`�����AYf=���r�|ݦM�^��L��0��#R/��*����oj��Vj����3c�2�l�w[+W�C{j��Y>v��욙�������l���}�n��YY�L?��灧����(��i���q����J�N3�6�r��A�A �+�8�!Q���vt��F�㊑ZQ�R��+NRq:h42��������t��R>@�c�"tQ��%�<;�2�RM���#��Rl]�y츑!Z����o����έ{�K�ee~�{�s�m��@AX��>�iX��,�\x> ��:wlìuF�D&��h�L&DT�$S/z%�����`)��S3p��})�3� 9"�Dz�1W2�0�)e��[.p�D�µ�b��X�QZ�m|؁pK+u2�e�-�j�����Z}nrrkk���[��k�+�];��� C���sL{����v�|Nm��?9>��G&���ƚ�R�MN��#h�0#�E������w &��$KQ��;V�
V���t�4ѫe5�R��</�	a'k�+�RcVC�%)�𷱿$>gԃcdIԝ�9v��,���<����@A�瓝Y/� �?�`��	�3�fT���E&,k\���sBNonX�h�1�@�a����)<��A �|��^{2���h6���Ɣj"Qq��;X9��0�&��M&�aÆ�O?��{c/5��a]W�8Ƌ>8�e3��TN��DjW&��Junz�����U_k�\���cn��导c1�*{��k�֤��k;����};�;���g-k6�[֛�sqGδ������R'�zr�Y�Z��7y�n�����1���*�#'��D���iH-����$,� �� �l�D�;����Aȴq�H���Ag�I6�:`��"���@eaN�EmW�Q[t'רC:��2�������v�(�Y���eT{>P��� L����'?9�6��N�pϨa� ��aϩg!;�͌���0�{�8^ ؊9����Fn�G����w�oQ��;�x�T����<��?�	�Q[R~�;�xE���eMxes����!�{��H�r+5R3U:ci��2ͦ�{VL�6�f�[��]��1kn��4�5䨿�D�����{w\���Ϙ��[1^n�N��J�VjW:�A^��,���8��	'��9�4^��R����j"|�۷��]�y>�0��D��J���غ�46Q0�h���,�`���t,�����Дy�A��=�fmٸ�Z,���ۿ=����]��g"K^�u�c��.�o�狃���<��|�8���\�B�a'ƬdQ�����`W䦀չ��kz��e<�4 L�.��zأm�u�V�G\5�g=��*:��qo~繹 <L�o8X���L�)C���}j1vd��k&t�&��67�sD��y��{D���.���Oz7�����p���So�;kd�4�\��j��i��>�N�vܳ~�����zm�?��/ݷ�وv�c/{׉+v=�S�������?eyj./��R�B��f.�xg"��Ĺ��t��Ǥ��>+���X.�fi,����H��ܔ+C�m�p ��  �Ah&=hPFm&���=o GM���T��I8��2�  ��"WL��F6�� t�I����l���΋�శ}8~�7x�g�,����3~����j.֐-F���ڪ� `eY7;�,� 4�5�19�Xr�m�\k!���>��e��c��q/z<�����(�T@�6����C���84D��I�e�<���LDr�����3�YP��>t��҄#I`��J�r�[���2nV�	�ҷKS��9�5=��o�?z��\��l�����4��������{�}I��/XU�?�֜��߲�I��zf�0��]&�0��t�G>�'$��Ս�8S<�9�L_7FL�.�/��Ĝ�ј�)���?��?�,���.ai�u��0�0����1�W����y�%�X�Łf1 ���C���!Vv�le>G����$.3e�! ,� 
�w�w�k��q�@X ��q�#�u���X^m,�v;�G�_�d� h��I{��/}i�&��	pрIlO�RJ�@�X&'m��<��B��2�,޹���t:��箾���<�IOZ�dµ[���vl}���C�0 �3�U�i�9���c���=�c;O\����E����Sˡ    IDATuO���g�����w���ܞ�k�Vfó��J-䈉�x�� �1I���K�v�ַ��uV;L�C��#s�7�1\:�
�$�"�������&��w�+殺�̘.���1�����}�p�ا��� v"ʮ����-/E���^*-ulb�&7Dͽ8��"G�Ar,2.�9)�"��f��d &�ꫯ��a�N8�	�_��_���ш����)��@��E�������ZFuv�.e/ًԦH��	�n�5��3�]2�'M��wd�`�Oo��Qn=������yQ��7(?��uѫ�F�\���͛_��'?y�bl�@\�L�����̊�U?�����w\���`�}Ҧ.�=p�oMn�����=O��'+�v֨����X*�K���Ǆ3�k¬�۽����.ơE�"�L��;'2��8�AV����a59�.$@�}��&���4��t�a,8@�$�u��`i� 1LV�N�*;n�$�����8�?G�T�81����O|"���Q��y��8]H@N&� s�pm[$��l��F�j!9�p#R<&b�4��T\%���s6��jχ'lzMm�� �a˖�3\���Nˀ�4!�'�F���d��U������?�R���96�E�V�}vÆ�}�S�z�blv�&|�^�~���1�Fy.'`o��Sg�q[��{�Gw�]s���z�m�)����+�����tѲ���c͙��R'5K�y&�E��?=99rX01���5BfE	�2{�����(�N�ڀ8��!�Æ��"󛱔�� 7 Lg�%"���Bg��$t@����7��ܗe� :PM�_��A�p�a�׏�.F������u5�{���|�DD `$��%�6_a+L�E��k-���Uc�vŤ��7֕2	�c[\C@D��w�7`��`�b��=J@�rp<�g>����lX��; �@F��,V�Nd�>�&#k
v�R���ƍ_w0@����c�s�p�6-k�֝��{�9q��z���nԇ_����ZsԶ��M�}׹��{l<�K�k����m��]��DG�Kt�**y�vޝ��|��&�F,S�9Y���@c������ʯ�J�<�){n?�:2\-:.�K�q��=0a�4sNx�X��v���\��\�t'6��	�vu9�b��R��b���������mʅ��>`	p�l�� `NbE��u�Ġa�F^l<&l���@*d5Rx��a#8�	'�'�&�]�;֏�� ��&�0���MS%�]=�kRâ#�?�  a����Rٖ��x>=Fۓ��n)R�0O�� ���/��u��~����Q��<uPm�+��Єg˕�_w����?;}�	��c�E���n1�{�M�NW�?�����w��̩V}Y�4����I���p��/��3���cn�@;;�Fvg09����d"֗s\ygG� l���ς�7,�侔A���PF:2�� V��z���5!G o8��/�����l����\������&lG��]����8]��O����*1ۈv��`��9`'��� ���Rmu���(��?+:�Sb$�ep���\ĳ�l�76�A�9S 4���3�F��`�7eP�Xj�� LY�YڌVN{��K6��L� ��\�n���l�0 ����]�nH����������2&x�
~�����۷^\�v�]�G�*�6S��]B]��4ӣN~T:��3�X���������ǚ�UG$؁U`$]ѭd('��e�'ٶ�`�%F���L��c�9	;����G�e�^G��xc7���J�e�Pf��06�}(�0H��8���a5�خ�\�Q�})�sr�:������N��8qE�Xǃ���; �$��cӡ�Wd
0�:� ��[̑A,9�n�),�KԌ��
���@Oe�����2p��;@��q��s�OAI��I�H�-A]����b�Z�qP�+��"gt��w��kq t,u��9�6p^E�W�s�R�37n|��1�Em���,�0�]�Zz`�q�O���n���_��Qz��9eӻ3q����ݵ�7�7gO�V�v��*�+�Jn�N:!��ſ��kci|l,5���j]]�����t؅Ҁ�vtB�	��N��g=+O�D�Mfg��}��N':�M]�T����ݡ�/���� 	�����$���;`QtD���#�-Ĳ�E���ܶ�2�DPv T�z?�C���	{ �� Y�20��F���E�=�A���u�Yy~ ;�z���xGdA�{l���2O��J̮I�)�ڪ��种aĬ�ע���I�r��B���Dw�(��+��Ю%/��mذ!/��_�lk��#y5�����O�9�x~�՚+�˟ްa�	�2L���X{��G�~n����o�C/�1������;Ϛ����V4�>�Rn�Z�.�M*�N'<��.��rs�T���z��#� ]���^0�=s�J��b3�Z��h)c��#G��e�E0.���_��.�!��+�`5,��ED��H�9l���ʈu�`HLb�"u��bp�]�]��n���^d\��@�+S�z!����ds�>�%�� f�2<!@�A�$P֫�>mړ6 �hK ���Cޠ]yw�Rcܱ=mM�<���x��F}p.�b����N,bC������g	��\��B
EG80�\�_~�<�>T2���y�	K�[�"��������=�3��=v�-��z�Rt��^�ɿ���[~k��[^����G�*�Z�=�J���d��M��	?rb:󬗤j��*$���f��r���KC���e��x���
`�A0J�2�	�+�As�	{� ���ɒ��눎�B�saU�J�ɽ`($����` �a��2E�Ƚ�Xb�/A��8�q�g�}��f�e8�m�Cu|�m H�h�<�̗�$܊�>�'[Vo'��m@���H7���w���Æ�x9�c[��@�bsM��͔���[@S2��|HD�@d��v�_<��7�$F9����IN��v��="�a�0w���;8�=�u.x+ō'��6dY%6�;�$�	\�1?�i��A�l�����+����@��91��y�c>=��Qn~��YhZ��'m�n����dٖ[/[37}R�2Smw�R���*>�7�H'������Zᩉ��nv'��v{>�A����LBi �u�d�z����,�
�-��he��	�z)�b�iuDϧ̰6�Z����T��6��(L�g��`��ι��cȖ�*?;�3�I��I��2���D�������$D� ~�^�=Wtw�`�\�kB,���"�]��U� );k ¬zd�מ�� °W��6x&�Źh�xI��sh�N'��=�kڦ*�I6԰9VJπ��EM�kEF���xuf�}��x�����xhw�8�����ڰa��L����}B��{����ǟt��xMw�C�z�5�Ԧo�q֪-��Κ�=?2V�)Ä�U�J*��S���ؓ�����Y�@�hu��;�C`��>2R*�	;Y�F+@�M\�'� G���9�s�F�� ���r��������\�9@�8Sadh��f�j{ ;��E|%�q}&��0�v�������E�+ھ��n`<�yœ�~aꌥ耰��;yw�F�$t��/�b �=�7���t�#���jK@��L�~͹N��,�/�2^刮u���|~���}D	�ߌv��&.�G�C�6�]{��0����b���mګ�Vh��W��a�]��kN�������M������~����7^ݲ����l�t���*ө1¥4Y���N>!�uΙ�����R��������D�B�U��#��QtⅲEw����7���_W>>׏�8~.��,�w9�spY��5�% LP?���� "�ᚬ,lqy�g&FW�]3"��@,��Eh�H*`����3��������, ��F$�����6n�-Ѿ�%>Äq�ѓiC�Y��xC�O.�0LM�g6O�A����,���n=em���>���q��'��O��T�2�~:L�L�v*��se����(Ca��1�uw�y����1�R3�aQkV�s����kl��c����~�c7������<���󸍟Z9���WOn���k�{���S�5��6Wf��&'��U�צg��ϤR��N:�Ĵlr*���lwC��H\��]��6�52B�#)�����t�x|�C�]+v��Y��;:'1���V�	���9�������6��� 9�DB����;�%>�%�ΚG�x8�0ug�u��8�s���۫V��N�2t�Q�G �� L�	_�"�ri�G�6�d�6�@�k��6��b�y��QF3�2������a���Mm�gs���c]x��z��uE�NC������hO��>�ܴS`��!����3����}n~��z	����ʭ7\�~��W�g�n���I����\J�j����c�g��������L%v};���n|��m[ߘ��e�S�z*7fR���J�R����������/����Dj�Y���E�*�a��
��#D�#��{a�t
2_ѱ�p�C/�r�O�C+Pv▉��;�0 Ё	Q�3"W�v��vG}��g�	����/oT�ڟ�^�sd[2E�ⲛ �v�	�c�|T�Q2�����I `r��	S ��O7��m3@��e���@ȵ����=��1��,,bGp�+��8pM�E��j�� '�%(�;.tr��fH@,>��y�������D!�C�0�h�K����
��6�'3E�"`�\�Z���_�t!jh�v\��	��@��Z�j�S�J�LuC��?:}Բ����,j��RT�3����*w�������dgv�T�����Tnv�7�6t���T�=�ݗ&''�o�Ư�����nTD���F�F��AX�(~�;'P����P���x̀����
H=D���Pnf�)�g���Â���0/_��R�C&���D��sd& <�	kqp;��;��j���y3���] 󐛁�u��~ G/	ǐw���c�##�g,�׊R��b�ݐ[�I��3���(_p'yv�KYB�r�w�Q;v~������}�h�E�1��z���Qtnq�2��ā��Bl���~Ll�T�@c�Z�N��Ax�ƍo\��7^�v��� <3τ��~�<��Ԗ��<��/׏>������~ ��s�����o��_��{ǅ�=;�9Ѯ�f=3aB�J�Z��ȧ\M��qg�Uӹ瞝�y�O�Nj�z�;����1�+���;��E ׵uFZ�HqcqAa����袟;� �Ɓ�c�0��U�ݠ'�iGaY���+��޸V8���; ���s�L��zǮ���A��G$t!2aT�`��?�Êڃ	S�)F�X�~�b�c9�,�XO��9�- ��}�ss��f��}��)�xM����jM��R� ��sb��A��#�0@�����e���}����"��������9�������3E���6����M�ް� <vˍ��ٶ��T�M�R+U��t�R%͕ʩ^kͭ\�O�cOx���1_��Mu����~��'/�}�'w�󋝙ݏK�4�棭z��]�N%�����t˖�R�\J/;���'��͹41�l> �  ��y��0�;@d�<"F�v�^d]	�h���^l'�W�2�8����K�,aP>�r�atb\�Q�4T���L���Cd�����!0���EX.@';Q��B˄s��b_���= as���xG ƞG�Y�����߂�e3l,��`ɮ/l �m�`	pAg��F�oT�+%6Wͩ�82Yȹ6�AqQ�����0��*):!�)N�.��/��{�֕OH4�8@��AC? ��c��{�ڻ�]�����N���V7�D�r'uj���Z��}ԉ�j�#�����q)*e�56m*�X{�s��|�-�����R�������ިݚaX0Ӫc���'�����87����f�����w�`x��4��|\DA��ȋ���p#iB�<���X`Gh Lg�?/u��ϻ��������bd�0�1�c��t5����3 �V8F�c�Ja�_�n��P��.�l@���o��
�r8����w�3��Q^�+�6��K|,@(�.L>��m�u5_�-F���W�qxs�.G(��<�9y��*�%�u�,�n/��A�Xy��+&�)3 N���R�0\l3 c�\����p@Y���i�Ub%�_�u��z��z?�L�+�n����۶]��5}T�<�zk�E���DoM�ԩ�ӞT�4W���1'�oj��?��i�൜�X�cN����s�+�����s{�����i�*��ޖ�r�������4��ؖ���ү��/�S~�������T��r�8p=�d#b"K�E�sa$�0l#f����0��lh��ha4*߹-����u�`	�8@P$J]�w���N�ŉ�~Unǖ���Z'/�R�	��9�C��d��T^B0���vڼy���/ �<Y�-��}�M�CzDX1vc��h�zbf5�q��=����a�������zl[%.]Xo��)#�xõ���ye����9 ��C<��;����q�xe�{��>Pd���6�&�LD䏃L|�Ŵ��F/�߽�D�����eC@��0�,�T� �ϲ;o�t����hͮ�g2��[ޭ���RJ�R'ͥj�WW�gc�1�8��{Ձmq?�2����o�8�z�֋V��E+ZӵJ��ʬSn��'���c���.u���8:�Fz�ǥ��n��f����Ra!�(3���� \ԋl@����߲#����1)��VL�=��8 j�"���� � �	#IP&�W4�Q@�q�Ƽ����c*up>L���fۑ������(�Q-h�HGqr�g��mڴ)�2���d¸� :� ��&�8��.S.z'�_��O�m�Uk~�{�.n��GD Ҵ#�y�l��[d�܇Հ���p��v��l`㑈p=nX���_"�������m�6('�}'!x,���(C�] s*�͛7�aɶ7z���;jj��oZ����Z՘>�S�)Gnj�rj |��4��33�������cW���\p�(F��c�������<�����wl��W5�{��TO9�|��:�	�%n/U���N'M��R�>�M��jtݤ6�]@Ɛ^��e����Fo'���0V/��wq�.v נ/��	�zq��� �!U�%h�<#:�0&A�c�dγ��I
�B��Aw�ו>��;���#�At.�lLP���>�腗���W�` ������h��!u�{n� ����Ł3���A5�Y�0n��,�d�X~���|t%\tã�CS�y��(\5ʻ�2�z0�D&\x�eH 1"����A62*Sv���>�<�F��\�h=t~��>pRe�7��s��Ww�M��Z�]�r�L��f��j*�}|���Tk;��]�͹G�'�=��;^��~^w]�7l��t�g�߽������_&K�&�i�!�d�x�>�l��Ff�,��Ɲ�q��1�9�>�H�+��ҹ�4�� �я�c�, �L�bXLܙ~���\����OC;�w�S�I�{�b�5v�CY���Z�r �&��:z4����;c�A�:�SP� laYx&HD֓��^H�_�3:VoF�6����w�!^#�Ɂ*��L�+tRz��XV �]H��9Q��F��
�Q��Y�{�6{�a���8���$[��/���x�ٜ��� N��%�����_���-7�κ�;^��5s<q©=;�0aA�=�J�r�-�Ӯ��={V��������>��k[�,����������2q����w�󧦧?ٜ��`���"W(;� ��w��<Jw�	�J7�%��l1�Wt��_�A0C��E�l)�1׈/��|3^��b����͡;6;	D�0 �s�j.�'���)2�����s2��[1Z�/����f��p2v�A���k�J�  �IDATtQ�!u����"��4�5f{��V�c�@l�5��kjkʆ 0�a둡GV�5�������`��s,:=K��đW /�d��=)c������%K����ౝ��^���m/\՜9�]�M�v=U�K��.WR�Y��N���s�D��k�jc����������f�66$�tC��M�R@v�"�&2J?ը��q*hq��GU�6?Z	!T�(M?�&�*�
��T�U�4���!�/0^���̽��9羳g��ݵw�����̽�|��9�y��u�4SH�^���]s���6�۾Y��\ɩ���_o럟8�.^xP�_��?����u��8���BKA �q�тf,;+��t�@|Ǫc$a�lȓDH�C1P� �������Z�� L�<���!#)��]k�׆.=�	�9b�G�y��#w ������Z�C��]�����[�TSDK��-��3��N	���#�7���I��[�:�A�.��~��F>(����o+�F~DŭF_�lJ ��?�j�C���<=|5�Cz�vp���P�����B	=8�SY��5�[3I��v���g���?�	�<cn��+[��=����:ώ6ϸ��P3Ƚ��6�`:����,��@��\ԛ�zN��ު���,����G�vKc�TV����f�>M\z�M|tW�^�� �c��u����C&)؂k
�v&o	[��XNF`R@��gu@�5�_��MGd���I�A���݈ &�x�� �6M� ���@���D-4R6�H4C�Ǯ~�^��	�A�a4B��$)�r4�$��E��o�k*�@G�^}�U����y�\k �A�W� �)@���I/�2�w�JI��m��,=P� o�7�s�<2r#�����>�.�G|	���0ʄ'���pA;F:=�oS��	!&�'���?ڷo��o�Z��Ov杧�?����3�^e�Yd����M�1%{�g�����3�gU�����~�7��w�wYe�_�rx6)�LM�p��or����1�llL�f���]��ӫ��z��LN�U����hvz4Lj�%�0$,��L'��T�I��'�� `��I���#�`R3I�؊��.�`�F�du�����#�L2�0|a����(Y��?���э�ɠh��&�FPG���b��cF9�� -� �>�`���/�0��� ��$y�-�݂W���n�s��'�A;��yi�`�A:a���6����3�`��Z�.�v�$�?��0<S���;T���qz9vA�3 c3�%�K�w-���������_�+��:K�0��d�G�qݹs��W����\$y�z`��;	$O�m�Hpɐ�A&��ix��sΦ�d�R)�a��
�t}���I9<���=�K1d����?���ĮQ��j�M�PZ�F�R�ګ5ZĪjU��Ԫ��R�����V5�ؔ�����γ�z�s�3]��p��i��L�0�zo�y)@TYfvf��LS"-zDm�0z�EJ�Ę�y0P^�3�����=s�C["	��sPD8#���ﾶ�|B�����o��'	w��
�	.�S�<r�qҟ!��&�Rf?i��	��\�Y�N�mO�	$v��ģ�bHj���qE�ʉX�T�($E~���8�kq��~��s��~��VǈQY0�<��wm�3n�*e(��!2Xp)W(^FYȏ�M���ڐ0z��(���1%��Zp�À&�N�[���U�rZ��1�Y-E����X�:�%����Aio��ޘc&��g�����w?Ek��8�-�6[����j�1����?6ٞjW+E��M��q�F�I�6���F2�����D�< ��D?��������+)��n8E�	*�������V�m*����2/��}���$Q�� �+!���6h�I�5?E,�qI�Ʊ�6�:e���� Ì䠀u.n(=�f.oZ�*��ڌ��tZ�O��.x�*uS�ʩdKҔx+��$��ðc����:�ԸK�,��M� \����5(��k����wh�l��h�m��"�Κ-�Sڱ/�G�,{}!����;�~���T]��q��\���o�X!rB�:A~AǮ�w�ґ~k�D�"%ᭉl�4Ց[�<����3�XGP���:��[<��|^�8;�0�&g�7�K��8��B�w�n���aEߝey>�o4��v��%��4D�e�~Ʊ��?Ӿ�CM�5y��w�k�3�����d��%�G�o�=d�;���I��<�G N���v��<������0n�S����'� j���"�C~�Ñϓ(�<�+m�z���{@I���pY��9�qʇ
�#��O|n!�}�T"[��*yy�Z3�g�f�
����<��>�!Y�CF�����&Gk�sX�yy-®����2vW?-�ʁ����g���,x/F0��H��"Ax�Qu�����?�R-��p[�<���1�\�Քۡn�G�f�d�%���{�𞙅aF i��qee��#7� ��3��׏7���;$��iX�z}:��`�����LuB��?���<��("���y_���[9��ED��\�P��Q_!H���I���B-���M�B3jf�={�F,�7j�I�6	)�8�_V����>[����wkZiͨ+D3#�0��0���o��?��y�Ʃ7����?�?�:�>_��~�����Wn�J$����-�y�w-�U�!7�=�K���62���U�f��7	���	��I|���*,-�\eF�I�G��Q��x�銃� ���}�tW�B�� я�<�.s�վԣZ0y;�pE1��±G]�x~�s��duF1�T7�N\P�����K*�d�5H5��{���៏�d'O>���͎���xr�&�{�կ�B�;]Iwȷ�*{���Nŭ? Ѧ�Y�6���5Ɩ���Z�g�n�M���d��������̈́�+���]�&Fܣ3��ȝ����\��m�����J%�7�N.V^���lOI�W`��Ԛ�;��rFM�hO��&kSkwK�F�d*�=���e�yU�2J�~��s�<�<�m$�ȁb��A����F�1$�JCzG�9�0�X��=@��L\j��nl�˓�7��d��4�̈́���=E@���Y�����Y_ވ�o��N?�vҖ#b	�
�{�� %�R�o�l��u�i3����7�( �0_#G����W:�z�F�I�Sh�_���Ĵ-k	y�E����uh|�wrn�I���K]���+ԥU)�~��J�M��h:��,���0XyO0a��W�m����m�	i[p��������b�w,wk�n�i���2���|Q�aӿcOd�����ޟܟaP[_�BV!�,��
���I��ʠ�5W� �>���O1*��T��C�".C��±�$��&�^�o,k���`>������b�=`"���r�ʼ�"���T����n��րj�����B�������!�������Ѧ���C����I�ǯ���>ZHc�K�V��
�;	�`"���X
���/�����$�Ďv,�[��5�8��f!�-F�[i^�G��b�#�ۣBb?B�/_ɋݭК�Gb��xI�ݩ+��@0Z0c��]X�)��"����lps�lU֩ʑV
�&,��焾��;�E��sx�g�k���=���qH��/z	B�=���@�!7l���������Y��K��WCNC]�����:�0�w��0����ɻ	�%�e�4��()��c��+iY��l!{8� �j���%�&�Z0��ә�<���Pf��36?�[�z0�M�?���x~[�੓I[*�" ���.�$z��Y��f!1����>�g���D��UgΔ��2%z_�ֹ�\
���82�~Mg�kTZo�%s1�ˑ������ݣNw-��)k1��o�Z�F&WК����D���i�5j��W���r�mEwm;�u�`��IP����P㕗~��Ka����B0�A�q&�>B.���0בTI4K�� �i�?�R��1u�03<ԏX�7�˂%'�mj�9h���^����ivJ��A�P�4R�m^���P�MݸY��� 	3�ܩ��^	���E1�5� ��$q��lJ�O_&64��%*�����b���G��O�w��;�����F8P��cfpBiN�-1R<0#-p"ϲ���R��,���a�F��IO�sd���e3����I�F�]&�N��74}$x{L��*۸9��ԃsNVق>����{6�k�9�2���[չ��y�0�H�e�UKGd�V�)��
�?�R�:���l���<XIZ����l�j����A�h���r�W��y�8�X�;��쎈~�)S�v�O!��ێ}. �B���t&�Y��)zG�A�2y�Ÿ�3y�`�
��PeuW��.�id�sĻ���r������!?j�6�#ي�V��}�;�v��#7� �eqe=��q-MgDbc�,����<�=��]79r˫2���x3�ȧP=���}���u#AQ+��|��CQ}�Qűq�E���Ȳ� V.Y`�F4���w��o��{@���x>��	t�@h��;KmO+K�ҷR+��6,.��+2c��A����-r	��Y�����WZ,c�����2�*���1ۤJp�����h�J�������Z@�8�/ILM�����W�#�'�����J�|����q��ٱtǀ���Ϸ9��wW�wB�B�lk?%���������Κ�ꨭ5 �_R�F��Ԯ}�3�"��'?�2�S�t���(>����Ν�O��\��p2Z����4h~{{��8Z>��#@�Πu�Π�S0�.���sF	Pԭ��d��H��=��PX��x�v��o9q���="�J��[P����{ǭ����;o���NՄ�6��.��mE�������Ҩ(���<�պ�?	~�W�-e-6.�$���ɋFaZZ���?Ǜ������cU���!r��鐵�����ʗ;^';0i9fI���i=XI��ɝ���:��^�\�n�{7��>Ԋk�����>�;��Z_���0�7(penHV�3�Sx:�Ҹo�<��{@A�4�t,r�A���hqb�&�au=��S��
��.��E!��;\�(l
R�Tݖ�V�^�h����Qt{J�~aulM1��Z�'�}��:��~ϝz���I��`�ϊ<O�.��GS�؜��i���{�k��	�;�j���\�Դڹ�,`��>}M�=;?֘����D�bZ��"��V�aH=��ov��,w�pn�ө�o�Q�+�/?$U䴐�^��g�:ںf�c�j��д^�w'2�_�&.F�m8�z=E�T��|�����^�*`���r��.H|):�F0�ޟ��_�2���2B;���P�D�	��3�'y̭]]CGmIR�����B�|v^�=�}	�߯��5��M}�XI���n���2�S��ToO����ޖ��_E����KPɸ����Im���ˊp���D�l�"G�,cC_���G���)��ui|ۯ�u4�Q@N��)j��3�7zœu
���hPۋ������|�q-#&�1E�vK��/j�ET
#���A멃�,*-^�!��GA��T*u�*��+�6�6PŁ���\e4�Ҕd���x益�������m��Bj"�7.��̗m71�!��U����;<��o�]�K˰�u������������񏯣�S��FB��tC�_WW/鳇Z_� Ps��k�Ѝ��x �����ö�nv@9��s.ƒ�d�������%��V�C"��Y��n�qX�6�G�?��n���$>�z�c��,� �WF�.��}1�{����
W�+g�VK�Kb��6����w:Z�%�Ko\(�[�s���������2��=��($T���.q��hB�@3%��]d��a~~GIɿ$�Y����������k�*�[?Ceg�3��rƔ2��v���ގTڵ`�M�oOl��PK   �yDY\��䓝 Wt /   images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.png�	4�k?��)�RB�SȔ�M��(B��"2g��ls�Hl�D�L;��"2�����d�f��:u�����}k}��ֱN�y�羯�w���~��sAI~�=�0�ֳgdT1��Y�N���O���j�~�;u�����*�{��-;���gͻ���w��jګY����cp8�uKs;�+���V���d�=�~�Y��#F�ͭ۩n��J�5ǆ]��_*^-	�w�s���b�_����v���O�oԽjV�kw&X�]g���_}��z�X�C��Cї�J��EBxU~?X�<q��8�][�����[Zvۿ��C:P�}`_���)�V�,i�)G몁�{k1Зs�-�9oo����׌�i'؅c���u�_���rO�������9�n�ž�#������HbgO��l4��7���N�/R�
�PSHJ�M�+j�g=Q}�O0���+�j��nvl� ���4�3E�w��|`K*�t/f�ש�P��n��p]C+{�QY`:o�|�'|�݉��	z�g�����vL�ݮ2�	�$��86ױ7�x���-mk��\���9��晭��`�~^Uj<K�7�?�Rw�8!��f����s�v��U��E]��,�Ε�m��O��]�7���:b��c)x<�L�Ѝ^083ٔW���;v�<]<RUL��8#\����IY��+o7����촷�!Nf�O�Ń���2U�7Y�9����?�O祣��R]�G�ǎX�6�\�O������BA:/U���1?�z��^D��ޛ���������\�A�:X�����e�}y2����}ǩ;�n���:ś���|��j
��.T5�Xv�@~y!l���z5��8.� �� cdC�q��m����F�3��F|p��(�tm�~� ?�(����A0>�^�<C��Q:�R��j�P�iN7W�����9}�n��8w,[ ��s�Uˎ����b'c�����l������s�8�>e����<�=��\Y��N������/���ԥ��j�ɚ����V5�螟�qF:&��t=;�3�%>_ �S�Ҝ��!;�6Mn��%3�;�=D+/ک��d�G��Ar2��v7��gځ��n�J����O혳h���4��&�ڲ�i��^�gj��z-��G��Kh����RH���ak硲9��
z9wM�Aj'��A��v"o�_�-�
1�m�}�����<Š���!$H��X��^���1�ZJ��T�I�m;��x6�~�c�5�����)QI:k?XS��RK�#��	Zu�0չjY�u�!*�Bn0v,\�1�5^����	)K2
Cx<�-�p�c��ˉ�	�4*Y1��E�e=���;U��`�h(��+c�f7�LI�{qB�ez_%l�²��"k��ǋ$̦Bٻ8��pt�P���M�#��Y�"w��1xYYr���� Hs��\Z���X�< Lu\pY� ,F�$�����Ǻ���<*���(�ZMUAY�hZ^��vB״�*lާ�����Mv�]��* w4�I��*�H�RG[�L�:��Y�QmY�J�s���gy��e���A3= @� �ϑ�#I���� 6�����S2)�i�8�ɧ챓��������y�^$���v#1u�vf�3w��(٢�l��,Y{�I�G�~���+���_��&5e��H���p `��k�k���E��v���H�V �~9`���Saq�?�q�l�2�总�>K�Aj��j�֭����d��M��u� �:2�:)��q/��H��	 	l *��?^���uލ�ݽ�:r�,�W�w�t$o��^�ޖւ��B.�#����<�V��zd��Mr!���M�H���wl�5�p��3:�k��-���W��M���룔-T*u�AfA#[ǳuz*��G6pw� "��j.�R��L�$6z�XyFuܱ�pg'w���:6�x��̾M=�����c[�7�r�\��S�,rW�Q1�A���K'Ɍ�\�l)�v٧ᵜ	(��s_p4��$�/iC��X��ZH�^m�{�QCt	�Oի���NS <�eb���ʸB�V�!Z�8!sp�6&<4$��BH_A_br4��������I��i�
�;���8��͈�ğ%ƾA�J
[�z�j$�7B��7�_�"Mf��nkӭ����ddd��4���ݝ���L9ONM�lٲE|��R�=<<,�R[�1���o�+,���������m~����\�v��CV���Q���"���6�<"�����!NΞ�G<�Ǐ�jL1��ٚ=��������E[��������������1 Y����+ Gz�E�<��;PE�)��ƙ��H�5��=z�С��b?�'vk��>>0���]�>`/��k��X�?I'S��]Ix/�_����h�꣌bL��e$�\�x��@�k$�q�s���v>�4!'^���n���F��@US���Eg�p�W�fA����go6�H�J� �9jq�4��fWm�� �k,aNԶ!�e������y�`���Z�$�%ͼ19���bt��3Uԡ1hРq@����Ψ�)�d�  ^���Al�Ν;k-3�8o>V�hN?H.�'gQ
�Eqs.��i��Ғ�p�jG�X��N�g���8U��\#	���KJz����9��;�#���@�E�TiY����U^�i8
y>�i�$/�����0���� I�PyzUM��	<��Fm�E���e��i;�S��cRl�bσ�Q�������8���6�|2*���ZQ�n�`�0l�����	,I��=y�M��3._�R�Ԍ=�g�^t9PXI������*�IYj�>��Ǖ�;M�;vݢ�Χ��<����`bbR]"�4�����c�)����)�ec���/�w<�%I���ݽ�dJq>�#��ґ�<�F���b���}'҉\�F�i|8Ŕ0!�C>�ȮZ��X������V������f(Ɏ��i�p\���ܭ��X���3�$g�BlF��D�.�jm;������H	�)
�W��DŇ��T�V�W�!	�F {7��t��6��f�8�-,�FHyH�6�\A$9�TL�u�ac� ����Di;=��Z!R�rc4 �G:v�\#jg�e�㎝	��6�<<.&������D�$y���#�/�)1�Z��f��J�$9o��t��h ��ǌ�sFFF��s�k3�\�@ �� #�$��jdO�#""LQ�=� ��b�g��ʹH2���>�TU�ep�J�� QwY�8�U���g����˙�R3���?�"3����X,Բ-�DH����	QQ�a+�-D�����A����qN����Xl8�k�'��E�9Ոv���3�m�D/�� ,xq���a�
�ny;�}Fss�L�ԒQ�4+������P�	܍��ϴv��b���}�I�xgr�%1+�R����nSBb�e	S��W�m�989Du�C�V�aB*v����[)�}<6�-Ķ݉�cccg>�0(**f��4��I���,͉�O� t�vѳ��J*X�J)���ik��>Y/�1HbZ��o)�*5u�j%Z)5C�����ȃr��z~)�S	�B���[A� P��2[=�h~܏������F�̍ёX��5#ښޫ5
��w�n0#F�|� ́��{�T��d`�eU� ~>��L��P�b�gڙ�kn_^���7ؔ���X~�Ƈ�\���T��-sVf��!W�:(ks>����q�d����¨ց�6[�fT�$17�j��W�;?=�+p�����g�n03���J4@�G�����v��� q>D������h}=:���,��;D���U��d �L��m�=F�ə�/�>����~x��3磹���[�NQڲ'�Y�&kIa�a1���*1��k�T���Q����6��=�,;J�E�N=~ <r��s�{|8#g� f�����!@R*�ut��/{��|�ȶS���g�<9�$#3��\���;5wy��K��~�B��Bv��x�N�����.O��&k��SV�zJ3[�u�j�=���Z]�,�ϫX�^a��<�:����v�I��Q=�Qu2_�b ���g�v��ܩF�\�fPɫ��F����'��ë����gff(�ε�E�l�"�`;�5�����&ȁ�� ��[�	t�9a�繓l�S^6XX8��X�W.miI7.ϴjϙ*�='~4����+ęS:F4��ɿ�ʽ0�㢢����;�O_$���I�ւGORKlrE�1����W���<˰WĲ�P{�rJVX絅S'�tA��	$d�ѐ�dAJ��8��I#I]�#n �n-�	�����$YC�L�\�~����e�8�u�#��ܟs�z����yd�'$�R���bm9k��*�E�.�i'���Ea[=�Y�
Q*��\�m����X��rFm�ER�:ݨ}J�
��B\����N������]J0�dF@^Z��<�ӵc��__�~Q����X�B�`cx�2�^<��	d!i���PNM����sʀ��^�l�)�.
K����x�%B9�i���@���D�Dzm\R�O���ag�e�>@CߩOCM�M�g����)����3y��m������G�{����s����0�4����h�
���G$%�
��T����ܜ���O:����Ú
ܒ���N�/
'���r��V����1��C1O�+� ��&v=	�{'M޺eKխ�:;��F'1ya�-[���&����ß��'�K�:q�s/]f�D�X��S�v�s~�\vr�|;%p�B�­7� ���m�O,���"�s�ԛ7o	�������+���4d�ڨ555fm�9�c��J�G��֯_�M��E�:^�vtϾ}����A��`7#�TF@Q��S����y���=�ss챗��o>�Nz�$�C'Ӳ����0�Ķ��-����m�z7._��@v)�#9�<kЪA<�B�Q �s">˅H&��L��e/q�؞�R�����p��T���$� 9����u�@�d��(2�5/Bsꌱ�:{�����4G'��ƹ�)]���)5{6n2œ8��"�m9Cj>�Jgj3��DvT�Z<��	n�'�l�[X�ȑ#ۣ���#]�o7�޻�O�c���(�S�|WWן ����ҖM��J�UEؐ����tۥ��l����0?������nU��r���A��,����F�\�u���Q?<��-q��ݻw?�j˪@Y��;���:sۓ��C��$��V�'���}O�h)����Y]���qJ~6o�����=)�Ao��,7�z3���2 A���[�:��Z�p��H�TEIy$��;U:�0	����d&n3��ff����
Od{&�2���98��`3s�J��K�y��U�.�H��͈�1���v�5:�����`�T�չ����mqP�ggԌ̖m� ׉o0�5Nr��gzק�����i<^;)��q�-l_�"��fc�8�N��M���)Ԑ�����gTK���(U�	n�aq��ԟ)U��.�����`������4�Q���aWb��+�J-x|ُJ:d��*`��kwp򕗗��m����Ec��<�iJ'���Q���'�Gӝ�l�+¢�I�V��Y�(��0��-W�g�fc_����Mg9�@����1���E�������i��6 .�����tcE����W!:���(��B�D@������k�=�w����#P�rM8yU�3.�|(b�YX*	u�)X��qC���>̯�s,G��FI�:��Dȉ��Q�ns:�=�:Y�l�O^�ڎ�����^���jh�w��A++�P�kj.�#nB��y;S^���d�"��D�x�GJ�I:Y��IU�>��`v\تc�ÇUB���)�=�����ŋ݀u���,P�(�d�$���\�/���1K��l-E �q� � ��l/�R�q�"���!��Z�>.�NP�v�j�����T�������SM mGZ�<P��8���S���l���M������FID8:5��p�2.Xlx��*�a��M��O��
�V�[� ���PԱ1�c��p �$��q&��q��&��h!���=���3�>dP������P#ܔ�0���Es��S���y' �I�\���.)�c224d��`-		G�}��Ճ"m7�a>\�f�cg	�bb-i�^|R�_-W$��3���Z:�ej�CV���Q1\��o4Wt�E��v��@��%��?�4�T��ͪN��-$$�cU]X(����I�� �������;�߁�Ѫ/{����og�E�=	�{z*�"y�`Uh�G<�66��mV [�9o\�b�>|x����aaZ��Qb��h�����@�F�+q3�E���lA���l����,�*�DG�bo��h���nŽ����J@U�>r�B�w����,�M=������7ɘ͡211]��]����Χ�%�Ǩ�L}����'j�|�II L����(���[��C������{{��zP��)��v����ph]��t?������e�� 	//o�ҁ� !�|����q�N&�?y�j �4�9��9h��a51솢�¤3�ŠY[�m�]?|�g�柵׊B�tr��X�U����h*��`��3�{q^P��R�k���Z�z�p�l��y���Z��r��pe�3,�����NV��)UT@C{�W	�R)cmED�O���Y=7撮�ˠ�A��K��j��e޽��6n�7h����	#�'��4Fv,i�4zm��&�j-�n�˩�,�Ï�B��\��ʌ����?{�������N@�px�ʝ1!�>}���=_������=�Ү��۶�'�����)���p�\'��I�P�	k��8�:5���E�ha!o�_F��{ �P����g�Z!�=E����l������\
�]�KӁ��������oߞ"���x����LLm)!�ϐ����}dT.t�c���:�� Z���M�n�v-~@�銥%?99�4O�����~ļ���(��)̈S����N{���hǉ8���� \T���/N�^��y�_�����nC��N�[�1��JК��J�� �w6_?�O�LF�?PO.����'��V��8%F��9>�1�Ɋ�B�pc�<(Z�rnٺ���ֽ��I�J^𖃠*#����C�ub�j/�������e�(����G%$X��yp��L�����f�Cx�8<��ӓG,�M��y��e/Ī�ܿĿ�dm{K��7@M�ww����p2{'y>���#���=d���Y j>�\��'���Ă�K��Ǐ�It�MT�i� �>�A`�i��[.��;� ��$���X8l�d#��SVUAPT�����iYY� 0-5�r�BuB� x8�j�n �QX$C���K o ٴ��+*+��f�Z��`I�����׎��?`����W��MR��+�~l̚�趶��!3���Y�] ;�N��ʼb$?��Ag�����Г��l��?�z�T_�F}�Oi��'�'�Ų�Qg��� F�}$���4;�d�SP���" �����Sw@z(F�O�<[�!qMH2@]�����0��ʣ�K�x8p��h�3��k�,}�rT*A��Y���w�\�_or����xb�J�B�� ��J?���k���Y����lL-Xt��FTpD�&׀tz�& ��'UQ�qh;�	h�JJ�@,YP<���s�ű��e�rvs��,Ǚ��T�����)x������}������������=���rg����3����G�3����;��D
b�U��	 ]!=�JH��7�������X3D� ��~8s7�cqH��J��!��`���a?�-$(#S���Ufk��F��ƭ-�S9']���i@\
@��I���9�)�f� ��-�B�)�.�� +�h'�|�ce��.�4�Z�=o��u)�!Z=�����kI��tx`Gyz�f�$�9�q��O��烍w����'<�"g��(t�~��bB`�K�Z!�f�eW+�6�,1f�H��c����l�\@�*�>���R�Н
$���T��J<�}�:�>M��##SV��a2�#�Y/%c�M���JW)6�b�t����=�^-���%D�"�»<@�j��}F!6]\�4�P�d�5�l@bdd�3�7�O<�r�HPsIU���"35��l><ߣǎ]���3+�Ft����H`%ϣ����Դ��[�c��r�m���PPa��S.���v��%t$]�#��[�faf0jm4.����x�A��̌����cj>WE��)@Z�]�b�r��1�j	�.z����+Ϡ#Ц4#�a�۵[�5s�ym���7+��V3�<PdT�;6�0���NP6�F�2�,���� g8ņښ�?��"2�r�ږjd�s��ʊr �#�� q�\#�\;����� �+�k5�h�`�f��B�'i�v+7L�]��P}gn�H����}�e�xG:����i����?f��`N���X�^sy@AP��d���*����0(�>1�A阮Q�د[��.��q���TP��H�gE*�A��@h�ĽF��{��2�'6T���]sV��*��~��H�0����NZ�;������U����2M����ΫW� ���p��.E�i5B+ְ]%4��T_i'�!�b��]7 (0���\>� �󮬟i�W��qi=g�E�^�q�F���( �!h�Y���$�\��O#E�*�̰>R�[74�@����r�Yf+|�~��E�C �֤��yތk�xߜa�*rګW�XxWO���?��Z�m���2�z!�;�ǀ��qD�$Q�%W�p��F5c\Y?��[�d�������YQwKWk��������Ⱥ�$w	���Yf�LV���gavR�m;�[>��"�'�ycw[���� =D�[x
Wn�ViH��y�Z�<��h^Y���/;4���V�R��E��I� @�>d�~9`坹�t^v�����::@����l�㡆�=Nx�{�V���r�Y��/5����-2j{�7h��=���x<����ͥ/� �,��m���	�M�����W�3�o]+�S�����m�Ė�I�I&�ϙ�m�D<�y�5�����(IO�����@ 'u
��r�	�+x����A8Y7{�P���~�=��+�3�B~ et#xǩ;T��qǔ���e�MPCt�|1p��"0��HS�ф�z�[U~���D̢�_���.?�l@*7���|��[1䩄�h��88QQ[�n���y�|*�c��XYEq��nP�	�|��w���9x�1Q
���H}�Q	���k��/--� 'N](x3�x'@>��UTTMN�C�"..�{��fl9��*ׇC#��vniYm��l��8y��zfz�)߇?�2��;A9�I����Lgq֞�E����-�/)u�BCC��9o���I�z��n�Kݞ�_�|�|
�?�7$�]�Az̺.]YX�X�<_'6�F�L ����<~q�B8���Ig�,�-`$ɨ�ŉ��iQJqq����@�؎��)Gq�����Ԗ���t^��րw��8�7Q��6��>MY��W�d$�[�8䦵[66��>w�ꞯ_�3�Zn�[~�߉����ǝ�:*L��?p���-��O�s����d�ۈl^�	�ݔF��	)�1��q7�*T�LdR\�B�wg����ygɊ�>HډH]�v��q�����N)@��b>�VM��y��F�q-��@͌|����UϠ&C���G1�����w�7�w�7�w�7�w�7�w�7�w�7�w�7�w�7�mÏ���+���_��/o葆�ʵ�o~F��|�ESV�V:o�XsH�=�t���B9�=�����6lHz�v�'�D����{~���)����=�v��RG��e��î�:{�]��f-�0��%;�����e��3%|�*��6K������"֦�A���A�+����f�g���҂mn����*)�`3|QPSW7�aq���B۲��͛�ʒ�k��y�-��L��v-jc0Vִ��Z���)uCA�	S�^��%�kfff���i���/߸r�GP@�bu]��]m�F̘��,	���-..�222.u*���,Y���^rñ����@���?._��[�YXl�{'���;�ܪa����*����H�pC���k������u�p��`���-~�V�,�I,v�oWHn�pȀ+4�"]����� �q}A���ۅ���i=��I����c��sh<�A�:�\����+k����=� �Hc��?Jv�����*����yt��n��
���ޖ�?lC	-�Ǯ	����v!(x؋��θ��(��R���:��NP��'~��!�`-&��L�$h��ӋU�;X�쾵���3g�A(��8va�)����N�/�@�O�%j ���2�޽�Qq�QK��1E���1���)��驩�SH�s}��2E��񟹛�j0S$H�x�Cg�V�����#R��d�z��d���L;�M����ۺ`���跉m�R9<�e��^�-ߡ�:i�4�?��4W��|5�A*�˸��K�?���rER��ݱ~c�*QUJ8S���ERػ�}��U���ޖ�G�M瘯�|�ʍ��y2��y�E��LV���#�����:u��I��ډ�i�s����EDJy���Y�QuC!�g�Wֽx=:�\�*�i��0I_�#	����V���o���5>_�81��p��4�!?�S��c9X��u�٦�������ee���l�2a��gN�="�i�Y�mF��ڪlV�b��}C|�;�9�A����J����zV�/A�/LM���&$�i.`�����]d}��%�k_tH� S�o�ݧ6�����eF�U��0�t��t�Mf�uq����l}rfh
v
.\w06C�~by����D����v!��.���ɭ���t��o�i��N�<r�R�d�6$"E?�ABfTf��ej��͸%H������KVD���<�)g@��lw֞�C��_������fi�0c��4s�)x1g�;��o|�O���ĝDov����F��]�Ѓ��>��Q`ő�lwמ�EWT����g�Z�����u��'{��y	���U�]=�؉�I��=�Hi�*=�I`�
4��]�=!��Hr���.Խ�5��5;����#-��� ����.��|K��\�dD�[�Ǝ��U���pڢ��0~n!]|9������}��D� bM$�]�G���=�=�^3�ۉ%��+�'sǻ-O��-6��߉�{8�b�h�9M��]���EȈ��D����ח���WO�hz_��-@�?�>5 �/���-7ڞ�R��A%����y��o�7�	��3��7[�}��^?|�e���H� �|��Yki'��E�_q�,��>L��Vi��AL��0k���y��h��?���|����0�Bj���Ō�Y����k�:�Өb���t�+6���aRR��h�G\��%���"=���;����ͪ?��޼yiO�݊��Ҋ�-��E�g6���f��C������փ�c�!z�d��5���bXc������׈Ý��	��M�F��d��gZ�)� �D����Gz���5��]w�A_���e�����b|�!$�n��Gi���U������Ⱦʚ|���n\�`?5�m�Y?�f-}��ҫ\S����]�(���[¿4�����ٴ�8�0!ˏ����CBC�/�V���-�@��_��Q��';��d��^N���$c�IM����AC/������Z�n����h�
�`�v}�|��zV�0�1Ӌ��O2�"X�/�o�j})X�=E�
�R�4Z�v �ێ t���[���������@�^xL����6�з!r=�� ��I���`?"��R~�،�@��yet��� 3WA��X��7��4���8�yZ!G��W'N{�ox��ߒ�#4
���l*.M瘪���E9�0�y�S{/,l�K�PU��>q�g7b�B뿒�K���Z,Ɠ�o�CƢ�v8����"�%^;��\HA���NV��8�E���U8�$la�^EP������Ѿa%$g����F�K��&4<��3���{I�`�����x�e{�
^>�-PN��nf� �E�����f������Bl�kKِ���Y�i03P���@+w�-ETr;�����C����"�}Z\(�'�S�*���|=�8���8��1�S0O-`#hm�C�h���2�=����<d�B ?@��˒��!Q����ьO����_��N"�3�xF��N@����]�8#J�!Ǽ��a��&u�M���&�a�,�ؽ���8����+���g�x(��� Z;��m_��ɰ�E�s���T�>�u��F��.�����z~ ��L��3#d7��������/XA$��?�lTc$s\t�B��뇂�
�����l@���މ��h6�l�H���,e_� �Hl���A�z�*.!�|<<<��
X�q�3�0<��^�%qY�u>�Ve�~ڪ$�Wۉ���z�w���-�MuD���pɏv`Yu;��x	E8k��)���?��N��X���'��m�-�ۉ0�4gUq<���	r�����3Uq��F1���� c ��X� ���ԵkSa �����;;����ݳ�0k��Sؾc�´c����V���D�����xy�N^�Ի�EZ��;㌔%O)�	��N7Y���oO�U����\G���߈Y��%�	�v�*lEl�?�GE><وa�H�����W��~R��R�3��B�z���$7����
�������9$$1�9CO��J9��k]� �~v{�b�4��f~�{x]��T�(�f�&z�����Ca��h�S����Ok�7F�Q���>'�a��������WT�e���2r;�b!08މ�æ�p�̨h�����V�x�O�ڦD�Q���׉��e--O �!E�B��h-72Q��w��/�Ϯ=�� �sV�y� �e��ˌ����ՙ�ӛzC)AW���I��Y�O�L������Y��.'���3}�YP�?�Z�ztz�-�S�ML6��h�_�n�c���c
�(��iw��%)����?�*6]�t�h2wЎ�f@�����=Ok=�@��9�ݿ�?��X0���I�'@?2����Մ�b2\�l���'���O�O*4Ґ̚���j 8�z����;C:�5\�+S^E;`� c�����#���]��=�v��5|�#�(���m(W�@x�0�R��1��5�݃/�Ճ,�֞�p��$>�as�#���7�%�a�n��^���/#	'M�ȯ�t�C;����͠
V���^ج��E����<���b�6L!݊�~�˵2W�����6H��gP�@&�M9-^T��F}�
]�	.@Nd��}Z��%��܄���Z��ap�@��)C!���1�q��YSQ��*��[��?�mï�����5'��(A�i�VYPq����0�xƷ]i��WǺ'�#���E%���S5u�G؊��k ��l꿭�_�����?�%t��Ŀ�s�Z��a����������I�r�e�X+x F��z?-���}���wԕ�cl�p/6����,�	�!��8�l;Q'�h��Qv�j���Uh����2��<�M���v&��	�;s ߒQO��X��j#7���]��U����0��wOm�4=�����`i���Y֟ T}�F�/����&�� b"�8Ү�7��X'����?�;*�0F����$����b�M����^���i�$u?@�+hs
���M���0䈍Ϗ?�	3F�[�rG}�����f�<o�iVmb�����THV�Wc�9��I�+�@�MB��&*r�aRqd��3�{�H���^$0r^~�p V*7k� 	�or\ʄ��O���?es{�6���e~������Ʒ��G��Nn��뿭�=N���n�\���?�٤4e�9�\c^p�4��y�8Ū��%c����Kg��ˋ��-��;�����Bl�O�+��E�?�(�O����7�����@�|����\���`���t�k�"��B�pƟ��iB�b`������b���wi�ؒ�=���ڵt�dt�=a�b,m�ձ���6� }��t�Q- �������~���y�ٲ�t�X�
�w����ٳU�� Ԍx�ڞ�Ϧ21�����_����+`S}��*���0y����ʀ�̝�B�1T�C�H+�<(�ߝ宸9z~jd��:\�tB��c3�"���#��9&HaY��:�,37�ߺ���;v��=	�;��J�F��Q�H��V
�8�@{NA�G�J��"U�]eF��� �?^��Y�� ���E�>����˔Y�B���������6=qP� ��]6e�Ώ���T}d�݅Q�/S9�IIg���i޻W�[��0�yi��^[�سe�����e�d 8���b��>��%�nZȁ:�6  1�v�,}"��s=�hž��J5rNt��Kq� ��\!��?����� dd�I�O�ā#�ոVW�݌��6}{Ȑ�$�e��&C�d��kDm�Rȝ���ϊ�
�������QUvU��j���9�
T�;f��Z.���nnn��6櫒[䴑@��^�Ƹ �4pgn�
�*�J`>ӟ�Js�2���8 �)��1��ᰧ�"ȶ��R9��d+�@m���&�����	
\hLq/�ٓ���������jO��P?u�T�SHE���0���g�LH��[�n��sQ��ޮ�l�u֪`(��gn [�Vо�Bp����DdJ4t�1�煫�2��L�3��pUm{��.2��H�2�X��M���c�<�'1����Z�'cPu8=0���ь�Ʒw�w��L�����	D0W���!�&��ڙ$u�V�+���N  U��z8�[�tm�H��H����'�ƨ%�x5��؄���w��F�B��X�m'�B(&>^��*���P���7����J����������m'��[?���^�D(��t@z_mq*B-�YW��,`����5f�@Z�G
SFRؐ@/!8�ʭ{���Gn�WK[��fڛ,$$w �菲1�cD�����������5U�^�O��3�/D������UоO��P����iW-��	��g-`��d�;�NgR;91��,D�7��@hѤR	��(_�籽ծ�����՝+�౐����[:��#<9���0��=��G|�?p<���A0���v�}e�����|�h�D\=�8�E:tv��i;��7��'s6dp�;��1M@݌a�c���\�y���L$ᔦ@c�3mV9q�1vA�M�I��X �"b�WD$#�oli���vҎ�
�R<�n����#t�	wa���C��g��cUrW=�����ݨQ��Z#��*�h��?��J`���Z�|k0��bW�L�'0M��o�<���/;��|�k��&N�E��e�_}��ĸe���\th���d�<B�R�2�!h#��85�� �!�WH��r�W�ov�`��=�Z^�A���hU��� >L�>ubK�x�/(��+��?�X=#C���~��������=�ʓ�r������{1����>�s�yT��DtЭ��r�>^;����q/�^ϔ�q��ؚ}��3��[SY�8������N
�0���:�!�3�ƽ���}��Wδ��c�a��,����=�&݄�ak�f�w� >����-��Tsɂg�j-�l|k�J�@�Cb����ɓ��❄Jx���w�}�o�s�؆�[K�33����I��T��!VV�Í)P'?=��U�h���!#��� `�i4,"��E:�ɓ��6'Ǟ���L�b�?��ŋ�����[oͳ�GO����cos	$ݲZ�B��|�.`X�������ۂ%�9O)�~������6��8G���$�V���5�T�����G���B?|8KO���=�m������������0����`́����I�:�t���-�^Γ\��'�A>GOh��x�����Bp������_s����Ir�&��;����߅��{�<���[J�u&u����@V��f�̈O�)++��8��K[�n��ӭ���q��^�V�B�!���ʁe�8hL�����S{��{������H�����2��NDXx��z�|����s����>���5��/V~���!�l�~����S��+]k�?�w%�+�	��(}��gbbb)(�P���6�����EG]]}n)+F>�lr��>��%��Y+�@x�Λ.h�a-Ɠ���,�Nd�d�-���]�1�|GD�f�>~��#���rc�A�ׯ�y���!���NNZ�K�����{�u��rT�>~T�f��2Y��(yU%Al�;9�Jo��v�1#����37AY�r7�Ÿ��8���A�+w��r���" ۜ䆸9BE�ǹ:?&��9�!NNcu��4j�B��wM
h�N��ᚐ��-���c��~�ߟ+d���z'|���'���=o��);�[@?�^l�A��n�<��S�R���n��Md��Sԗg�{2�浓q*GCoGw-+))�O?Qu��ө���ߪ�㪳�����a\������!��t�ik�3Ǜ7����(rssy���B����(�JJer�տTs񨬪z�Գ�q�����Ruz�p������e��_0Hi4vw�gdd�z��IF&&c77�	�A�������_AZ�-,�~2�iΰ��:�#�ֈ$���x��~�x��T�^���hj2���P*��(`�)g����%��� ��?0 vt�PXD���C�)Gu�8�c�i0�Y�vi�7�n�A^[m(���?����DDD��3L���:?d�VCJ��t���cg���V�E
弲r9������\J���@_כ���g:�m�w�^��k1��e?մMdh_.��aqqq���f���#�CC�O�ͽ�8a'WE�r�)�\���
Vr(13��R=e�F��d�G�,��a��O|S�kOP2�Z�V�<�Nk�K[5�\v�Ƕ�ՃuJiP̦[�s3�t��L-BnEۉ�~��U��+�\LoF�T��@���/hFJ����x��������#Y%��A&~�{���KcC���Ѧ&;yUu�;�gf�NQ�O�g�n��M�.����F%TTW��d�k1��`�-����'<����ɹ��E��1��_r�q�Q+w�[.��E݌R!����=����$2�ZU�T 
a�∦3��2	�6��O�32:)�v��M2T^��Z�q��~���=�u�i�����`v3�c䲚2;��^�0���C��S��]O���
iY?R܉]9R�>H���8�A���S��E����/M*��<e�U��jZ��ϻ���S���{{+���Z:�����t}ӌ�`�L��i�z�ܦMOOW-�9�r��o�����LM��l�n��3
n���B�Y}���gز�c$g5٦m�w�>k%�H#E���>
}t�!ź��lfƣv`0/~��$��ݖ�b�E�:�Dzgj����z2Z���<`ဖ�~�ݓj���@�C��~>����C;(Ox>���<��R�A��������5��c����W�l�>_�I4g�G�3���{ߌ����CQr�E��B����V)��ۂy��p�H@扐t���H�N2���d��d�I�*:h�i��_�й�%;�a-<+&d���O����o
�ٚ�\�:Q)��B��I���޶l;�Ź���O.&4T�i��c��W.]w'��#�E����>(��\x�2�P+��.�	[(�Ap �������-o���P��ȳi;�t4������om��n��k��c9y0%����G%-����\�
Ni]<��A]���e[�� ֩%Q>��:t)��u�o�	ռ��(��
ְ�����Ns�ܝ/Y�Em{�y�*ɺ��@Q�wE��X�s>/�Ͽ#k�D��r�hc�ƶ��i���\OV:�ݧ��2C��]�2��i���i����a�|~~~^���N��Zv�����!����8��y�����;kY�k�jѿ�P��ᱥtH8M�aX��w��$��!A�б�7�����+`�/ �S�'Ӳ}SG��������_��w���N6 �W� ��Z-�^k�AҸN5h|���3���bf&+�:��8Q�q��TT��]䧪	S�b��J����5��i����=*"�	��7H����%%����A��c}����>+fRqɎ�1ݞ5��/5�e���`C�*R z3lv�{$�Fm�O]y��)��)s
��{�����'�u��W�p���rK2$^/�
.�i�+Sާ﷐��2�Ӗ�ҝ��$�w^,��D��^����W�2�0�k�H% ��?5�R��,'�t��,4��p�޿M������{ )�]��BY�d�*�@BH<(�9��f6̤*H�|j�Ce�Y��(�Nj�Q���{���a՞x}1%���hK%�^y�u/��@��H�ר�h~՜+�uJe��,��v����	NB֜p����3�(��7fW9����zí
�cq�ҹ����䅅힝�	�	�|��1���E��SEZ��)�̳c��Dvy�����.ԫFF1�[b�l�v�sS�G�X���5��W}�	a�VK?9�hU��$��@���@Su`,�4����M~�x|�k�@_��IƉh�u�O@�$9wƲ#�[MM��/m!�	��Y���7�҇�dd3���qcע-�8��7�����΍��Uy$��wz(w�@�VB�x��ͪ�g�����fy?ub�t� ��s�ý��S�aE��+h�w�\nll�KH)x`�q�%�P���#�.GiJt8
�Qr_�6%G�3Qh�V�#���$	9�PIr��1C�c��`0��{T[�����w���Ƕ����~�����z�.(u�|ك��)�/�NW	 k��6J��c������w=A�p�cgQ�U.���ݦ{_�;M��^-��](w}v@S.�"j�M%��� �`��Z��e���ʣb��9R���7�����������p�F	���LM݀��]�v1p�l'��2��( ���A�«��6	#�X��|����s@�+�33o���6zs�-�}_nn��'�ꩾJwU����u�ӣ�O�6�9qh�t_���(��<hmG+��d��M��8 �����6����W��$́���A��3�L��~`�+n#Ң��M7��@z�5�e��$�C�������kc9;[=_/�*�j�<(��lS@��|�v��A�я )$0Z�P���]��`�+))��5��n����� U����-?6�*5K�%����h�Wy�T�N|�� ������^rT�U�#T����Jo����_��Mml��&h͕�X�o'�X-�\����/_*�G3?3Q��SHD�F������s]�
��P=&�S�f�r�=�Z�_�1���վ�S�U��!��ʀ�9 N��C{�*�X|��2��p稽�x��ɳN>�\Nb܆������s!�W57���>
b[��yKPHzbH��+������=7��|��5`X1 >F���MuP@�.���0nM��ﺲ0)�24�_jȝ>EQ��wt�{0���±��Փk3�Ï�65�ݱ2�$i�'�F�������f�ʙQa&��� �~�^���q��O��?�H���R�P,W����|4/'⩒�(�j ��=o��-�9��K�@�W�
L���dq+��E�� Xt�$RH�<@��Kq�Æ<3��&����8�י��ك�"IӼ��}�+E@��=3����f��/'� �a;����S�����c�`i?���w3`��w����Ɩ���A(��P��
��p���>?�ذu��##e��������r@�
����C�W,�%�x��l�~X�oɅ�)�ߞ{p��U�#���"�� �e�,����<ܫ�>�M��i�'�r�q ����K�wJ���k�������4��jK=�>��m�)��o����jeB�G|,�����i���������LDc��
�z���H��*�l`��V�Kh���t�m�&�[�����j���a����r�\ ��QSS3�ճrF�^�~;�Wd��C�7>P�[�6Ƅ7��c�<����=��O?�pKꮟfHi�� F�{����3쵑�7�����
���Lܟ�|�;��U���&�������֮!��ݳ�.�B��%����^By+!!Q=�)ǒ:�h��X)�N�gx�yۯF�y3�^�OD��l�׽������ӿu� �?Nr]������G_&���%M��H���W�E�%��W�ߚo�l_F�f��p	)r��<�	�nj�u�'I'癙��/m�z����YJ_����+��l�F�����ࠇK: �U��"+'e"�p$4� ����h�j%���6*}*�kf��;s�V������|������q�������ٶ���{)�Ç���e�t���T���.�~���w� NIx��F��<j�������&����/:;?�v*m�w�fk[�f�����U����j77��t~�� 9��q|P#.��0��e�}����/��������W㱎��D��� ��y���U����:�����~[�0Q�NA�rV���#4����l"��^VF�dd��k��W��VY\,a�Z\�����s���蘘Ѐ� ѥA�(I�jC�հ}Y���{hٍ=.̖�$F'߱���Y�N�Dۣ!�Î�NrO�(������v��YϞUG��3��qp0m�RF�B-����r,i�V�����â���Ϲ> �����팭���0 �����������Ǫ������w����u�u�PKo����Zb����q]������+�n�9D��;s�� "�	 ���k&c�OI0 3�]d�X�q���U��Qᵈ���
~`x! �)��������@�ƾ�X�x@Z@ԓ��I|	�c�I��
9Q2�E~G���g��#^u�]F>�$"��P�l;Xn[+oy��q�V)��"��M�v���N ^��v����\��?�Л�ivdۙVB~^p���LY�l݅7��ͽY�L�@�����^���Bc�7R"8�\��� �^��W,-U�c�ΐ��<-~�ղfN������Q�RȶǲWwӪ���/f��>Tv�(QWW�E�b�W� �󯶯����i��a6k��+�I�f��WW+���-et�U?~�1��c����_��-����q�3O�:����7�����g�эc'����2�xڟ��e} Wn��V,O�[����c����˹�?��8�>��`��� ��b0\[�:-/�;Hs����={��i�=>L\!j�{LLL`s}� ��8{��[CY��|�.�7e[��vv>��Ѐ�G��T��X�}Tϼi/U�5������vM�B���n��IHJ��1uu���z ��8��x`��L�ĥ�=??�{�g���*������� ����u����8G~��[ /�����"��j���%���S���VJ���N��/�yzYK⪪�p>��^3ccO���۫fffՓ��%�;��۫��ҕ�Խ�[Y��o@��q�e	�]�|4����D��/#���6�����Z a�06�{��nLxF��i�������������ΤaC�E��e�nF�;�Ӧ�1zT|��9 ���\7h}|�� ��RލM����7w`jzz�@?�x��$L }O�>%-��"&�Knt]$YBL��u9~��U΋{XYYP��=����&`d��/"��I��	`�?���}�����nf[He��o���F`+Ma+v� ��]px<>Ɉ���K�<B�q`X0��#-��i��뽯|�����e�&l�����d��W#nm��Ow���ǹ����9��PW�(T[������֓��6�Ү��'mO�ʁ�- {hc�+��ve=}��*T`����{5lb�����^+ݓ�[Tص�R+�\�4��s)���h$�3��V�(U*�����E^ɫ%!'c��e je�;4���C�+�h��w�mV���>cu��D[�qkMg:�K���j�������g���_�4����8w�!N�oh�144�n�[��+s7 xP�V��6�Z�Dx�Т`Э�T�r�i����t�z��w|~��s��iƌ7;y�4�6u�0whge);=ee踻�5թ�8
���ި�+�v��U����a�k���a����i�\���=,?��0^����������vO԰��U�a��b`-�l��*��~������M8j���}�ڭ��%P�ζ>�mQ�& }\	윜����҈���"	;00���6�'V�b\Y�L7�u����$Rg�`ЋY.�_nW��g	zYՉ
>������믬?�_H=z��kȱ?�v�0p�K�12-�r��{\��QT(�`DS�N,l�O�Uz�<�C�'��g`[ȏ���jD����]�=1��E�C��U�ʬ��A�m�J�°�2I[�.Q�5��+���Ñ�? ��P�tiZ�i~��V"�K�֩gX~X*�X`3U��1C'��Wג��5��h3��_ɢ����V������x�����$t��A-֌�a�����:t�q1���2$�4�����A_Ӕ�l7Tϵ�4� �r����T�Z#I�� ��n���-'8QJ�����m�f��y �I<��m����zY�IF�@����~᳿H�L*���-�HG {?��~Z�Ն�
�2�3���)�7��"z��T1ޅ�CC!?mF�R����V()B""����.J���`��{ŁJ�J6^����M�~�n��b�/\�<T,���bfb��άI��.l��jj��l��j�&H]GҧG��1xY.)�+W<��"H������4���f��"��A��?Wn+d-�(fM[�{��.�\�25�f�E��Ti���������8�y,�@�Mx�$f�+ɈjЍ37_����bkR5>��u��m��<�
�";V��}�x���
�*�����@{�0�W�]y�c�ka�����
��bك��e��Z(�H^��;�8��ڍ�{�H�XL_mp����Kֹ���0"L�7��>6`��w|�͋��[+zc��C^����T�?v7��j�7����}�ƨ:�c�j� �܇�&~�#�*=���n������,�����s+�d���C6�u��T��<����߃�9�Z�C����{�>��.v{ &H-��+_��I#-�e����]��؈x���'�n=�<��x�^��сw^�/��b���T��4�.p4�M��ivv�����v�e]��i�&������l޿,8###�H��Hٿ[�� ��vw�y�.N��d�m�l����'"��m�D��ӳ���2A���`�&\MQn��u�����ۍt�ID�`���$���o�Y��~�����@���7.�FE�5=Uɝٰ�9�{e����N�V�4�b4Џ�9=�-�-������C�~�L���Aph�'��@�N��S��aO۟Ys�̙iXu���N�Q9�i������Y�1����x�ǚa咣c��������[��b������8�<f>���?�\¤=��/ޔ�
�����J�����W2�0Ң�:m�ߩ�����K9����?5$�U��>�E%%OK��I-�x�3,��6��mؖ����O� ��2h��T�2"����8�~����c��hn�%_��A�Ic�H2R��po	߳�Y��V֋��xds\��ZΕ�Aع�EM�y;�k ��-pѾ�G��+�����KkFA����xGx�J�c�Q����p�G����]�i�Tv�%�N��ی|�B���=W/��œb�(�߂o�e��wl��b���<�g� \q����S~ʖ[���d���3��cr2��Z�0�}V��YO�֙���O��ˢۄ,ye%��:�__��m/u��-�?��v�"+֒94�+�6Ҁo� [*�n��Z�	@�@�J��ه�R��.���S�!Qu�����������W�7??�1�-.�Yي����nR��9%mR6z����L�)��-�H��+���;"���q+՚~D^(��7߇)en�ҍOP��>����[x5Y�:�'2�.25��.��m��#wX��;�bE��0�5�&�#�*��N�.��.��5:.��;�蘹q�!w�G���7�L*s��>١�2�iԐ,-�4Y�f(���`օ�w�~ȵ��q�3Sv����;<����2K�{�:�Gh�&j�)h�����U�@�D����h{��s8C��Ʉ��&?B�K�dr|���q�ȵ5�������mx��һr#�{�k�;X�@�iv��f�����������]�Ƅ0�jc�:��z���*:�A���@~��ʱ�ӵޭ�홗��t�����f�<�+��щ��%m�G��$bJEn�U���a0ڼYj(V����T�r3���22��&ƲH+퉬s�@/ll��}.+�N�9��&*���&�<���ɂ=��V)_/��tқ��^fH
Zn:�W*B�`����7d�7�٠��;/\�ȐŶ�r~>�>߽�ǆǟ�n���`V!��[E�z��U��h��Htt��
Q�i�a�3��8BtdQQ�0zV5�1@��B��n��f~!��0|g�p[I�R��<�_9� b�BF�7��1�ӗ������c8$�0�E�t����=��mV��X��vޏ�ͲME-����ЧvX;�^D >m}s�m+����#�ye���T]n�Y�y�b�Lk%-Vu\�a�s��^��p.wp�'8��8aQ�K�1Q)��NS�0���O�踐���Q���h{�2�g��#�k��0��xهk���^)U'��ϯ5[*'�����ʣ�<�{��>�هߢ�G���P��g�>�Y��%s$�c)yB���Ǘ�8q}\	 �{"EY�Q]�(��#pw�_���@��6��K�ei��O�6����+X�e�_ȯ�!z�7��UQxݨ��c�7Û�en�<Zx�e�Y�ph(C�����D�N�&�3n�f�րi���o���!ħz�ge�`dԈ*}���'�>�݀�sK�$��m�uy����NΎm��y�>,��Wceee��_�d���\:�ٶ-95u�b�n�	I�+��iӍ��}�\3�;�ofN����l{3�D�Tٰy����ƀ�nG�$�ȓ�`�����o2G��_�y��{�_�ٔ	o����{)_O��L�ԌN4`y����u�/8S>��!�I�i�'���܀��:�VC�*%W9?p�7�gwҡ쒐q�\O�0�/��X¬�^�Y x����Ì�̹+]��������I.7��
�	����+.*��"��~HkqX��,7� �`�n����=Oڬ@����'��D���p��� ����c5���l͢R�V��S�*�Dzκ{�g&�������q=+횻��2A��;f�jO���	^.�+�2Z��}��E��)��G+%7�_v_�A-����{�����i���6l(ߢ&B�T��@�U~v�nZ��		'~���E!���5a6R�w#s@ڇ�]��1ap3�N^Xp���6B������*՞��:::��*��ܹ��[�X��;�^�E� �^����k!&-�|eHA��!h�X��ʫU��)cn�&�`$��퐻rԅ�MI|?Ha���2I��eц3���K����!}�O����0F�	��H+8H�,u�������b�sA}��Y����m�L���8�0��.����>����c�lJ��'�O���	=~���V�Y�|s�Z���;Xμ��9P;� �:^��n��l��͛7�����V�<V*ɩ�!�@rE(r���6�Ti@,=WC+oۣ��=�E,�/�~ɪekWQ �]��[���q6~	HE���tV�_m=9��p����L{��r�^� eq�9ϑ�bCa5��<��,6�lGe�Uj�{�XY�}y���$��=����jӵ��g��2���Η��Ne���f����nΐ%u1}�j죩��(�@�*݊��;��ک�
�(��s�0,���?�}�(�=��D<6Rn�aP���㉚���C�u�z��;�o��H�����M/.&v��i�����e����⟯8��+ 8/gBj��W $��:(F��.��=��:���|�%�T�ϟˋ�����#�CYv��z��)���6O^�
���0G��`���FG� �G*Nͪ��wX8q��V0�ޱ݃�ʈ�|y��Ju�H�G+pMdv�u��H�Si*�2/���2��=�o�^�?bo_��D���n��+��nQ��Ω���\��.=�Ep�C ��dF/4$i�~f�� vrDffT����������i�ϱ>|a�P3ݰF�N����{�Hn�I�7*�p(g��/�����l�n�F�X�oϟ?�02b�I����#Ms�N1}4���w�[8lk�<V���@�-�O��;.��U�����, �;JJJL��^���O[5]G��w�����(����������=�tD�H���nU&ˢS_7�G3�\r"�^��y<ձ���4Y�L)������!w���g��b�C��e�~\�0	�������>-�K��-F_ �+Q/���樫ѽ�F�׌�����A<=zT�h���prМہ=����q�.�F�<^����T���	�39�L[SЪ���^Wn�VSq�V+u�k�?:j�^�q��x׉0=�X̌�ޔ��N�xw4�%�	
�YEq���E�u�[.8%b0�CZv*5�f���R���||,o�*<edQ����ճ�.&\܌6���h�0r+SA��ڊ��V�O�y�}�?<��w~#�����s�*�"��h�=�VQ�X:�����PKK���Z0Z���jx�t�!M㴛8�0�g�koވO���u\4r�fld�>���Z��P.=��ߡ�ߚ�i쩪��
���G�役9���p�I��펜����(���"�圁�9���ۦ>��T�4t>Џ��_!�;T���X�f4=x��`��U������#!�(:�@'��"_�ǣ����|�M��b��JQ7S����5�(�� ��*�E����w'�����G�3�6�"�!>��#��<[�w��;�+J?��M��@�r�S⨧Ib����u闊���P����
�B�Ǣ�bG�� E��iSx[�ا�Ҕ�\�>G���䭘=&�^���+�b֎����
�>����JZRR�*{!!����_��!U�m��(�_��=9���q���� �k�~�^�Fss@T.����k��*��@u��k `��m,첤�X��^�r��+Q]��0��lt˩\,�>�}Db�$�ƛw�o�	� ;���uU���#zyVf���Z�e����	��t��4VzW��gn ��fKhM��t�)s���zXI��D ��P�x&�ު���+��dȢ���Z�S��<�5� �t�=��?���$\����R)7wd�tJ�ˬ�)�;U�mD��1���ۭ�W�룻j/:�[������CIT���Z>�Ϫ,j�c��M�܆P���+��Wn?����Db:K�Yy����Q�&�f�R�N��{�A�ǯ���!o�0�����@|�;���[��d2d�X�d6ڡ��q�����Q�^�&�q���<nP��-�����ĸ�].6�ژ!��˽�+���W.2��p�\&�ٜ���W=qV=�A�y~ }y�(]=i������k� 6�[��'�+��#a,�i��1�*���
�zU��PF����FA¼��4Z>�q��C�z"Cb��7�Q!��.�Zǅo��PUU��;�z�8K�q���9+��l��^psJ]���R�dB�UV���+�PG$��b���|[5�����O4�}v7�oQ��1)����?;SO�27���ӿ!�v�,Q/�u=�຾�I�QPH�)�����Ԭ%�LX~U��ϐ�S�"�o�Uy�F]Y&U�V�#�s�:�����ڬ�ʖ�� �=� ���P�G�z�b��e���?��o�lq�h7O�(�=�Ͱ���R��M�ڕ�d��I����С�Vi����8C�	.�W���SA��A�������G�v�"E�(�/v�+��pm��ۃ��M�J䌌�bcÊKn���Q���lRO&��$s/��L���VA��w���r�ƒ;���4�ϟ/�f�sgwT��8�����8ӌ�<$z(w8�m�]&��m�J��莠���3/7���4�WJ���kp疏8L�Eܳ�L+pd1�rA�.����ͨ�Y��'�7͇d��/KE,ݸ*��Z)d�)��MGG+�h������شo���Y�����1AY�����Ύ�u`�|F�k�!ON7`^�J�Ga��TC
K\�8{&�6"�[HĐ�l�jȦ�i���}0���n�I���+e�R;gg�~��Ѯ&�)༓�qZ����x�AF�D b*w�</�cr����|�L��<w�t��]�8��'i���=�Ya,��z(�r��x�R���:�
�^.&�l�Ϧ��3g�<4�a��^�|��޼�Wc���0�ԉ�)Ms�N����Z �7�[�ܽ��M**
��4&8k�.�L�`�aq\Pǁ逭��o�_9��fl~^�1Da�(�^GUu޲������D۵;������@�uB�'l]�����'�֑���fn��bΈ4��5L���w�Eov���^9YYM���������8~��X�-7rG�w�[��%8�T������A�����6�C���nd�W;�r �W��٬sY��_�KɲV��bHP���ԥ!�n��n&�[���Oϣ��I'�=�\ִ��
ك��.,���K@c�>KNUTT��݊0���´j�V+L7}�r��~L�߯!��1u��Ծ����%������d�v8
ݡr!]�� �:rL|8^ˎj��l%���� T�)dz~�mO�G>���S��ǸQ�&����<��	�#�(����SIR o��;h\����b�}r7C]nKU��a�����t����:n��
B�!�XK�@�͟B��,[q�P��3�v��*���L��X��Du&K��lrH�wG&��#�o��]���t���'�k�F�v|=��b?9�o�0�"�>��k+���**���D��Lfۦ�q��rn4���$��[��/!mmہ�|5��� �\N�B���������f�%Cc)�.O��yXT$e�̌��g�k�%��*���;�El��k���#��A vʄ�����MT���R�j*�VBb˅�vK��)=L�=υ�%s�|&~�lOdsd`/A}?-eU�v�gqH�� ~⢢��D>�������i
8��һ� ����rcGly���!�Թ�[}A�\?U�	"�Q w�����As������6g<�-+�����>;S�lB�6�S�����y(U��;.�m��W���8y*D�qM���X���ť���D�����^������ �O��9|�]�����S-P��ϡ�J:c�)&=x3^4�t�*��oq��Nĉs0��]�O��ݝ UgT#>�O����G�����̚<7K7��Ik�B�4���B�'2X0�j����z����>�4"��'
��^�#"�/����X��b|^��d+P|�ŋݟ�uw�b�6�S}�2��?s�V� ���!�"�}��ޒ����KE�<߀o@��yx�l��k{�5xR�c	Z.6Ѷ�'��鱸����7 S�f�mo0�#zY^`[�%��)h9ڏ���/����ע�K���O��hT��>��B������;�ԗ4W*j,G���?W d��`�H��Cst^-�������S[{5��q��9�+�ֆ>�X�����8��Ư������MLLJEx�.��������f�	Qt��7��b
��j~!(�����`<�tz��"$�d��fD������[����%ee����P�lbM¶�ē��p��gk�[��|		��Ç{K9I ;Ҍ���B�߽�f��R�O����͟?'�8��ݒoz^،|�n�:�I��a�4}�H
Z
>$`fZI�_�,N)�8�f.����֭c�ma�Ʀ�7�GF����ó�I��'�Y恂-Trꮷb�����6�~��,��H���_x<6kh+�kե���o�y�&��8���t�7���?�0���+A��� ���\����@�����(������+d���+����(�OK�[����<_f��� ���W۟�2rJ̗>0�$J�����@o9�Q��;jz����"����D�*�cW�+M���m6�:��Z��R@���������z"��`l�L��Y|�9*Xn/P��gn�G���<ϸbSO䉓'���-�v���ܰ�?ַ~?>g�8𨷶����d�/��� W�jb����������b� �Z�>¶X��f}���;s]��̺�!<�:r͙��~����Z����
�vS���>��	�!��3330cL�%kq̙��6C�������x���Ѱy�zu�x�����I�s1F3yZ��
�ZM-Gю�����fTdbC�5��h93���ϕ�5-7�b�㮌����U��������Ji�dhW�7i���r����ap���&����cR��}X�*z7�>tpy!<s\��ł~�a�I��H���
a���-�cd5��Bjd�cЕ�6�u�۰(J.*9'��v��_mo����FX�s�˖�#�+>k��n�a�P��#�� O/�<ŹHr��:��H�	&	7�� ���g <L��N7n<�3�A����5�S�Q=��3�&9��Ϙ�1g������/ͰK�)��$����y}4��ڼnT�e�A�&�^n��-NC2/vwW�^GG�x#��a�)a���}E�Y�a����O�GZFa�jt5�&����S*N��S�N�v�|� �@�����8���/�������]rGY���:T����]\9��kkR�,���߽��nH�Cr����c��W�C�����n�����:N̹��W�Dϵ�o��]��CNT�.�# +��� *��v���d��&:D2�c �r�6�WgF�
t�
M&=9{P\��(�RS��^<qQMDt���@8��s�q����͏D���2O�ډV��˺�5>:z,�2��^#����	�ߐ��'�x����X�a�w��.��:HnZ�Bm�ݑ���9����#UFC��wz��368��ZZ�v��b���%j����/pU��e���}�2	L����)�c�$����O��O�G(�`a:!|'SW˳u�S��%Nz�r!� �����w�HB��\�x�0�	�(��\A�����W��湐�kQ�˿l��J�x��_m��r҆��l��D���_Q�z�щ=T�!��5�c��&�I�q��7�x�pQ٨�D}*�iҙq%Ǫ�sg����۬$b��8��9��݄Z���u=�J�˗o�'�>\訂���$�;��'L����i�-\�,uö_\��Z�����
q.:�d��i��Dp� ��W�)Zfðm� ����C��_��I�jb|�==����rpL�w^�.|X/K�_|'Y��ȁ�4z��&�m`�ͨ�ɟ�%�
�2*6����qh��<�����E[
�ֱۆ�����v��TnOA��F��Efcf���	�������5�8W���]揦�c�`��R�~���M%�)�I���`9V+^�E�<�����J۞gR��<��g@����t4���5�N�[�������� -���ߟ4���y�A�œo6[Vr9P��.#<��3RX�L�E�7k��`�C��5��I%����t:�G7p��_1��X�P�������9�/���zB t>�~��A#j������ƋO�&�������"�$b���Z�9����Es�u32A;�)� �vªr��'���)��А����+���֗j_�My^=�	M��r�)Nk��
�*���+q ��V.��/�u���wA#)��!�9X&�~qqH�ԑSW��l!���.&P8(B���8��<Gw�_ǁ�
)C�t�k�?�;��7]>X$��:b1��oi0đ�I߄o4���o/Ӱ��!��#d��!-8Q���������)�ev1��~Ր��"J�[V�x��E��4���bOsg�U��뚕8�E�8Ҳ���p���XB�J����ţ��q�?�ú(Z-`��8tnK���&��G���mf_�.ĩ�}��@��m��P����r�L�lkD}�%g�}�C�_�VR%'��^+��7���n[���	�p��;�M��D���g֯�*Ӏ��ߓsz��n��`�<?��éqhP+�{k�A�_�Prf��%�T��|�l����GLu ���D�����ى.�HػYF8��!�h����R=�'�(�A�b�4J�5~vK;����;H�&�|����bcS��<Ǹ��i&�,S<��fxbe|��#����#�p��씦��ێ�1��X������������C�:IAS4�>��O���h��
��N�_��~c�ܤ�e�"�e*d��� y��#�o���U�B)����`�óS$q#����v�x��Ls��h���[86�0133���>���I�y��tHd�3��L<uIޅ���d�ȗ�촣W?l)q�������p��{���1�p8KS��#��V�b��[���t O���!h��Fs%��(
������a�s����EU��� E�ݻg|&��밸�I*�C{©�e��leVK�����K�=ٌ��x4������jW�w�ͅ��&A�J��ٻ��^�cklld��e��uSv����Q���7�^a�w�g`ڵ�H���8�8�S
gz�{e`���.���/A�e�o����h`��sku\���ZT���~YO\NNN
�,Ox��NC��u7r�(����r���9/H� �������wboųQ%�.�ة���
��h���P��#3sK��Q@�}:, 8���۴8;���e!n�S�v6���s3i۷��&M> n�[�D��}��[H��J\_Sa�_�؎\A���=��s���sr&k�}9�P�/���}.���cR��ܑ��"��	V�@��(��l5��5��CW��������V�:�l� )aӭg/�����-W����+0���n1Q[�ES[�9�u��E��������J����dl�u\l��z y�Y�ؽ{���L�E�����?�,a4�̝�#|0|n��6m�H��^|�R��4mȾ�>��V#�~jJ l*w�X��ڣ�y-���]vU�`��)������	*��ʕ+�0��"{Y~>_������7'Ͽn�L�E\l���0>��q�C[6f�5B�@x�_� [�qϿb��{@*jp�cWُ���#�fv~i�#�H ���w�G�*�&T��6�6,��3E�c���6X���ci����-��/Hv��>�s�%3�;]z_�=���E��yß��p��[�}5����K���K�k�`�9�_�aC\
 �t�Vea(^[ ���a�$<֑9�5,29P���7�a��`�훫�a{�U΍VA�F�=�m�|�����K+��?��U�5���V_ m��͛;3Z��� @��ȑx����(z�\�B��t<�%�z�iWp����<���z�|���E�����z�`^�B�V=bg2�C0���KDc5�]b(�cO�%m qy��KE`?[�����}�Fdς77�y[��Bxy+&����X� X�Z384�����oag��IK�Z�lׁC#�g�SkD�b�Kf���d�026��f3p�
Ѝ9%蟕e��7x���W��EM��Z�"L�JlA�\ZUޟV����)�8����j_El=������+0�8#΀�G9aB��'�4Di�PW�#g��{�z��3�~�Jfv��"�ɘ_�d���x7M�`a��>l�$J���6.-�hjj6}�5ð�S�:���)R:
#�u~'w$�dPKK����d���ߖ��*�<������N�������ͩ�m����:NS��OWi~9�j`y�k^Gc�qZ�z��c�B|-��̻9z���kg����s��TCNe����}���;�§zN@~�tY/�ꏀ� )b��8�H�.�<�|�1"���"�}�O��	3��{���/�X��5��Jj��2�ߘ�����y�1��S~l,�����������u���m7y�����S��I��Z5�6^�Gs����'+s��Zr7V��͉;�P�l�T���4�\���'3�i�VqqlWf�M�xbGǆ�@��T��1��o��˿�,f��as9v�_�5.���w2�I?��1� t�N�oэ�?���1�[�X��2��-JT���>:��z������9��˚�菮�?����;��Wް�����a����g�2���\-���.���p\�V�n�$_+誱��X1�����=nT�����E�;��:�އ�~���/HI�,��:��!��M˽�����<�!�<Z��g�\
����<�>��k��-�#f�݇aE2�s�k��L���	;�p�m_�9�ȹ�70Ӳ�;0�e��\�B�����x���1�%;���܁�4Ԥn�����^��n���6z�<��w�R%K���/�ֵ��*l��Gr>9��I8I�19yXSKK�q�`���/�q�ǝg���v��+ny̼ś�P%=����3 *��TV��������}zWa����6�:����9r�v��u9�o ��V(���ے��쒯wsE�U�������� 3{��N.���zi��;��/m�r>����-�9цԢ-O��&�W�c�^���7q1�>�(���^��!�g)~~�<�j�����YEXp��o�>�un�����&��H"'2�GJ*����c�o}�+`f7)���E��ξ��WV��/��� 
�5~S�o��|݃�c�MRڬNc���e�r�/��*��ψ���������mA�)n��p�]+�
_�=��E���k�jh�l��nO��(tW��9cnh8{L�0�:�C
o��Q��:2`�W�d�^ݓ��8Y�ᮞ�e`�%�mv�{�U>�)6��gΜ���e}8nk-r�{9;e�in�րɓ���>$o�s��^��d	pL�j!|@FI_�E���$eF� ~K�,%��B"K������aԂ_���c@���xHa<V�4c����� �+}{��������[�`uE[N�3�8M�"�=5�6o��*���o��7!J.����4>�w8������Sss��m�u]�H��qf��N[v��&�^ۢw�t%@&>9�y6뜥�����O��6���v#^I����T��#k��h;m�-�e��N���!���y���wㄶU�&" �#���̈�P��&~��q w�K-❿d8�\��n����0n����\�ᜨ���\���p-,�VN����S[�<���~��_pv�+�4��e���:�r��F�x��o��m.�m�I���k�y-xQ!�l�w����*g��f�0����-�CG�2?�-�������6��h!�:��| ���wB�y�c�.G�ݿ�P����e��{�ȟ���x.�C��ۻ�Ŏ��GI}��(����9&|��ѱ�)Į�u��m���t~׭�.O�څ������h�Tn�󔁯�F�j�5-v�Bil�����E�'o��4��%��cJk�*�=�@ݱ�Q���5�b�fz�͑��׾xj��0�R��F����r�[���]��p�oӑ����՚����xt۱���V��P<j�
�eJ�Ѿ�Щ����w@���,Yq�T�T؋s )-=qU"����>������:�rY�Ŗ��
�tQiZ���#�c���I x0%$�@ ���Q��^�rx/����Jn�X�Ѱ6��{�Ě�� ��ν�lI�'5�ڠ�*m��*-;�ǵ��������BD'C>��xx���:��Q���-�5���
��ߌVw�Uh;
�����P7u "���t��Z| 5���T��r��1U#c+����]��ŀ�֙�����Q��G��%}�ݏ\��T܎ak��J�������o��m�.�Z���&A7	�-k�&����1lB:.�pP�Օ������^�cgO������i�Rٵ4��e[�q��o�8�$�̾��2����co���.4��JwP�&��}wٻ��n�C�?�H|/WqD���f�'F넉'^��K��ߚ�@�(�r3џ���+9�M����q�«煋��;�����.?m��'\F߿b7}"R��6�E׀��C^��<�eq4ovxv��iH����C��PM��@��x���yzB������*�ae��VóR����®u�xi����.��ͪ�+��~�tQV���Q���zF>��9�y��ύ+6�}���!I�Z*��=Z���S\Io��Ž�֥���Z��ŗǜ�xH(�,h��Z,�6���L�d�=��TU����e�w���=��	G%%J����2��Z����@=999�*6��Y<c�>�'��n��j�Y��?.0�c��j�3�bl3��R���e��r�S��5I4ѓO}��M��et1e�
��ȕI�4�Ȝ���:9��$w&b.�,PQ���'������Rx|��#�� �[�G��E��!8 ��w�<Q�&&&���_N�=z��q�ؕa�݂w�ф3�# <��������y�>diĻ�^��kIl*�j�I�(��ڼy�3.'�^5�?k0�ie��pI*����p��q#�%��<
�B޽����qE�y�+��p��7W�&��[�>`˟�K�tM]��W��uX���CW��N˔�#є�C��o·��>���ͯ��|E�B�sx�/(6y_Zw� �w���Ʊ	o ��J����@T_W��#�~���\q���j��=M��?�)	v��"�b��&V�z@׹�-�@���N��hlR�ք���>�gZ�C����X�D�&�uVT(��9ο�Da��j����*�rO������h3��6��;s����w�8w�Ū̡ՠ���#��W7�5�D�"�U�����Es����X/����L�lC����6��?����Z��h�"����cI��E�"%�PS!����JYCҐ"I��LL�d�(f&�I�L��������=����5���6��s�����{��֥����=�H}�
��X�9/H�c�Ќ���X�
���:yg2����TeM2 ����]���S���T�,Ղ�]��M\�6���Me���X��s>�N�Y48�������W`i6���*b�>�g�$�իW�4L��8jXέ:�1R3J��"���CL�ID���[�z�a[�x�V�x@y��j8�t75��٬Ȱ_�N����G��1s���lmuuC�@ \�uZ~��HAS�r�q�i_i�K�/��8v��W'�GG�LI{:6{�ѵX����~6r�J���̞G�,�S�Ģ�	M���H<<h�*/'��]��������s�<<�=�Ōv��ݮ��^��v=�嫹ZBJve�if9t�C�T���.���t�����ڇ���]sc�:=2������ʿ�f剗����)K�Or-Mj�䂞xL��oow��.�<��J����eVcB��T��*=�hB���C�V�����=�CM�fSD�_NJ��n�j�op�Ӣa��Q�"�m@C��/�v�J�_� d� UO4i�85�5>V�A� �g�m����䖼wwŬ�䅺7�kF��5*���9@�]ųK�8���r��!W׫�bb3�ݗ��Uߨ���`!FJ��X����=r��$�U��1NU��ï׬9-�@?������a����I��ɟ@@��Iu �O�J �F�~b)����{fk�^��"����� ;+qڊAoUӛ�&B�g��+ct*�q�w[n���.𥛫�&x�< ^9��9̢���]������t�l���n}�8�h��s��CiՈV��%a͈�/[e/���9��tL��K/��P�ʢ򀠅�f�m�m
�H�p����[C$��}�:s��KVf����Mh&��c\������:z�hS�
��	n4���_�v�ӻ	��~44׊���j�=��V�z�J1�
��� iD��4�,�V��V�z�<v�)�K7�����F�*��7���c�-���M
Ǔ����(K�mxj��Gu�3� �f)^�e}���F�^�]2��Ke�g���B��Dk�Cmګ��#��Q'�=s��i�Y�h��w>b$9J�#�.,���8�Ǒf��B̊0�"�1+]ă��4BU6�t\���b7l���a��|;�Z��:Ds�zM?"i����#�m�Lz�y���}k�+�E��
r(`S������#�-��ہ��q�2f̵bBІ)� �̸LG��GFP~�=?�pu��j����a� ��W�;�!���z�	ү&���{������C�QR=�]�X���^���5� 2M|-Q���e�TGS)�Vg��Aظ~��}Ĉ+������-�c���˙t�f�,kL��ʵ̱�6y��?Bbv����GY߾�j����nZ�f@��}=��Ͻ	�zFb�ɢ�x\�������~l�g�~�������6!o��	����;��`f2���6�^����mR�#��Z|N��Ɇ����O�V���ܞu�F4���#_��G���D�B�q؟�ɛ.��7X7\��DOx��G޹_J��>̻�"b�R���\D?�M�4���9�?���^��RY:7�S/T���Ѣ�K!����)�+��H���߯v��B�
�Ŝ��)[P=Aдx擘�j�����[Ue������<f�g]��W�tH�%f�o�}iՍ&�|{�;��Kx��%��Ӕ2>�ۂ�����ĂD<OJek}
��1g�*^u��U;D$& N9>
5sƿa��$4��f=j�7���Z��ƹ��&�v#���j,"�G��̆����4�q���\���y��N��ӯ��X���ǋ�Ta���B��'�$[�N)�68xkЯɌ�\�]p�>��P�9��б5��Pd��a���=ڎ�&���"O�u;F��K���a/�9��$���/G/�f�n*)�ŕVˊ}�E��@�L��[��ľ�8�)����)�P��"�*Yqyl$@^��Ԃ�@u)����ɰ]��_4�E5�(~ͫ^@��jKs|V��l��jR�qc�ڟ;���6x4i���K�ىY��:���Q�@�������wr}O*2�Z66���M@������iuS��,h5	�	�w��뱧H�×������ϒ�wI���o�CZ3�K7�3^(Ԫ/���0� e��$��ԾֹXL�o��E�d����א 2�[)=�bq�X�z^IQfX&�uN=�#Z�mob�������C��.��3�c����\~��?rgliү;c iHO�Å���,�	���kϓE�a~@�X5�O�lY�.�(���sq�ۯ��ƿ?A4��t��|�ʑ��ʋ�0֫�7c��Ⲵѻx�滗E:�>�ɷ#aV@=�իF,:*��E%����´b,ŀ��7 �m�R�g�/5ڑ��I��G�[W��+W�L������Q �}�U���$B{2ᕇ�������x�=.��_�B�`�fu�h������%O8\ߗr[��{Ys����R����h�-z��E��[#�m
����5�`�(5i��vx|��0� ��X��g�o�G(��8��^�v i���;/�Ib|=�.��_׹0���q�w7JQ�q2���op>�S	#~RZ�%���\!��̳��|ݕ��!�c�G5�?@�e�:�W<�ϲ:Ӵ��p�U�O���e3o1r�T-�x�1�e��X}�T��ٙ�K�D��+h���̒HלK:��GT��߻��Ϙk���@gh��gdSm�U�B���a�!����ҢZ�[����:=�:�(I	�Vב�~���^��P���H"|����N�H�g��J��e���r�v�?5&���[-c��3O�_.G�?[��T�;nU��_6�pę�ݚ>�Xo�ܻ�CY��1ڤ��G���!=���́�Aʪ���Bm��;�����&/;�n��W0/p���&q�(Ȑptf��;�Ȝ176m�7���5c �Z��i�˖��YEfW��=_��y�Vm�S1���JvCz�Q�Rй��@`I�dP�)/K��rhiSss"l_%[�߇��6!�D��rx_%��J23�v��٢�Ǯ Byj�7��C�����ۀ!:r�ht+��r���2rx�=*�&7���*����bV�+?�(zdO ���jJ�#-%9�������b�)t�Q=F���uy<���C��#�Jgq��!�� �h��+�Z[��ȉ�-���8N�[u#u��A��N`�d���߽�!��g���muJ8�z�pְ�iKXl��y,��[�7�k��x"�����C�1��x���Uӑ� ��́��'�C�AT�\/�����b��-�YR��\�vlх ��#�IU:>����k ��9<��ʡ�3ԦY����^��a�Z���%��e������`���ʯBy�%S@h�d�b�G����	�iZ� aS{-�r"�-^���K��0Z�q��6!�h���7�ᗗ{5ěoT����Gd�_�����f��G��#��w�XI�!kW.A,���~��b���y�V��Y����w�a�g��v�;#�&4�e'p��]@/�.��	8a�;.�M�<K����(`K#I���I�1!ku�H@���߭���Kû�}�.�m\v<i��َb���SH��H�!�`��!ݥ[$)�k;8��ꃭ�r<.���E�NȉqYmN�+�x!">�U�j+.�}7����b}5����y�����l���ϡ_�ɏ�B�鎯VS@��tw㯥�z���TR��Aj���vh����Pql�t��B��ҹ�&H((��R�W2�R����98�owE��w�dԵ�@���h�b��E����ں���Z �����N�����W��Ș����L�BF"A�0j�v~2R֯�;������+�c�����|& ��CķY*���f_���/G�Q��J��1oJ�$P����ש����)b��� �z2u�~t׭�rk����U���_)V`:�#���%�(#5���'Hպ^g�?�y�v�R���o_8��b��3{ϼ�'�տ�'�L(���#[<�i�G�(\Ucj�J��Z�;���՜�v[�jƫ�?z���[R-X̀���l�)y�tV�j��,��
�Y��Ԫ��N1V>��9\�6@�����Z�
�;HF7�5T�q^���6^�ϙ�遂֟Z7���-�Q&J�+����K�w���8�X��}�T�?���tw���OĔ�����ϔ��*�./��T�v�t��z�tl��n���;Cb�]��[}YR\wC��*V���1ƯJ���r+mΰ6��n�������h$�z*YՄ���ܩڵORX.�'�V�?5l�
~aƫ�.����k)�L�˻���F	1k��=ǌ�i���SQHd��T��Ș��e_o&v����ŝ�M�N�-V*�[�=t��]�w�ZL�i��$�U��D��؉���S6�
��ߍ��+v������vK��i�VP4� �q��7u3�ƻ��l�����䞬�B�bp�k�˓�����K.<񖖒]-(]�U_��TavD}��|����aj��~�Ѻ�	�?�����N%�n�N̺x��>iw8��{���F�9�p�c�22V���t�'�'��H�����Y.�ŋj���v����{?��	�7������$E�S�-��嶺^�M�M�
"�#��i֣�]��Q\���B*����u�ۥ��U���Ք>�(��!�T���WR�z�a:��B
�
w�u1w���`�	�t�	��(�"E�&���m&���;�#Υ$1���L,��*&F����ݼ�rs=˺�!�����y2�-�-0�mw�?����uA��<�?�4���]pz��I��y'�1~���y�s����ս�a�%{=1t�Bb!8Y��#�n��
h�g��GO,_d��y�+;)�X��6\�����O+�8� ������%��>���*�,��J�e��g�Nt\U����V+��r8�qx~���߶g��,��b��{t�W�NɄ =,3�~��[+�Z�j�)&�9�2G ��ˬKA�����	={%�]G�?,�rM���7�P*��^���?u{��형q��T���s�ݾ�
��Q&�;|���A�̨p0�f�0�mB����x7<6�� R���(�3D�~�����B�ѣV��j�~8�����B��,�Y��b���x/�w6������i ��KM#��бF��L/S\u��W�s�*B@U�����r�i��`	%�& IK��2vY5������չ �/*%F���`����̜u���	
.�r�R���hK���+T(:� �S�����||+���NLU�9F+d
1���.�W�%߮��������%�!t���fAS-�q�|������J&-�N;�m)~[,�o�^��5{��pjD:�р�>]��~��3�����¶<y���H���J�\>)�(��r��OT�v�a��L-�jOv���'��3��ź{�'�wDsk ����k����u�K�3�l�y����V,���J�d���Ƶ��W7Z�`�5�������0-8�M��܆�S��>3$�v+�W���$��O�3\�t��������[����~
ǻ��W���y�[�k�b�oɾ�d��nh�;٫ =Q�u"сou��+�t��f��J���P ��.8k���nu������^A�8>X�z�ńr�����h���_�{_̼�cb>!~]�oG4-��%�'Dq��1P� �5#�Jh5�!�9���==lAȔ�i��� �z[�,��Ru��_�ɻ�p�3�c��f�\O]!,o�e_,H�8HC��}=�eI���0��|�Nu�1T)���ӭm��IQ��۽d_��h
ba8�a�D��dlh�� ���R$;��5�d�e�:h�Z?�-�˼�0�a����9m$�w�c���k���+��̓hM���?�D&ֽ�M{{��}�u��c���['jÖ1��?�������
�Q�{�����6,�&|{���3Ͻ���:Tҩ��Ru)�}�����i�R�L��<Sr?{*�35�'~o��g��p6<�����& ֛�JN@�)�_�t�Y?��>��9B	i�#4��~�j@L���R�g°q�N���e��,$hfv�`k�POЗ+|�>z�:�X�b�jg���(�f�8+q�����f�Ǵt��4�)��Lc�9�i�ًS�zN�Zr2w���|���v�����r��[ ��o�R�v[џq��ϊ>��R\Vq�נ��Ƀ�yv�,���$@�AP���������:�_+<�S�^oŋ�m�}R���7g$%��"u��7?uV���s�B�^7�`M0�]��B��I�{�A�k����?^�[�`�B)��^.�=g��x�?��"`���n鬼0�p�ú�*Z;�B���%8[`12��T?*�fǷu�l@�3v��5��6-���A��(�'�bJoV�b�ё f��;����T��a)[JW� ���ȳ�+3�
�BUW'���.��vo���\,@㽉�&۳r���ߞ.�����ޏ�������}�����Ѽ)���<N�I�R�a����ODb�Qx۩��e��b���%�nbCNu+������=8;,��s�T��3�M쮆�fc�7�()Q�������&�LdT�v@��6�WN�/gT@O �F��*�L'ԉ{���M��]�ő�{�Q�'��D��9v�K?��J*�_�d�B�s)��L����X|�N]j��\�c�P�/���ć$?�~��$A4�Dw�ϯ;��� �J���;^u�Eפ���5�X�;�	M��`l�*$PW�ށ�)r���ѣ�٬���
V�@ >D�J,<�	�:*���@6��f��o�Y�fo���,W6��Y��i�z2��z�q����3����E�">��<�03�ڦ�HmhQwE�;�>*t)�w:WD��:�ǧ��g��?�y�y��~���� 6.�����~�Tk��(J�*���ʧZ�Z6S%M���eB*	�Tq[�?ҁ���r��Xቬ��-7�d"&�qo"���=���**�O��su��ź}�z�B�����cCo�����Q��9#��������:��M|<=e�R�t%&ȇ[����W������K}W#�J( ���;�O�?�!��ղ���1@3goS�6�e��;kW�} �I��ZЩ8�?� ��V}�|�R?�(U�I�+�t�:'a�AiV�^i�ڏ�PIg�cjn-��/VWڥK�ﬥ��o&6����$���t�<e~�^a
��ct0���k�h#P'�%��|�h����GN������_,2�{��
eK�
��$_�n_l�{�f�ы��+��t�cg�m��s�%{��"�1���=�~+o7�s��G �!�D�g,]�{X������6k����O12�Զ~���ș}~; �ӄ�������� ��t�?h���� �Ж~9oxf��Y��?�f߃�w���s��_"��FJ(F~�Α=w}`ک6��P���©�����a �#{:�?t�D|�r��q}�s ���:�����y�B"���.x��zdb�$`� �B�*]�mj~�����ν��Łe�{�kQ�]L�����z����CtP(��Qh��;#!o�������ڝ~w��������h�lP��]��/3L�� ��ܧ��ԹS�]Z|.E�6��a~�e�����]�ɋ䲣�B?]���8�+vbJ�Gݿ?	�� ���,$	9vK��6N����b���������]5��^M����
�����@����ҝ5H`q5#�^eXؾ	���Ӥ�Ö&e�un�����j��4���),u=W�.x��o��{�k0h�(�� mH!1�֕��Y�J̐�Ke�j�|0o���B�
<��e�'�e+v#�&�H�E1�Hd�Lt{����b�vHe�q����N�j��wR���k�LXMB�h'��N13���?��=M�V� �v��0���z^�
��%�ˡ�h_tힸ�Y%˟��Ɏ:��1�A��!P:R������8�C�M3v��y6�駚��8��n�!�U���Hc�ͥ��Z��À�C
�?��w�Ub�z���#O����G�٫��{���i-E�]�K�`NO�} ��T�����=�~��q���e|y
�%����z"ӟ�!#wBO}��-�ȤIcJ��!���S ���b5r��ߍ��Hg��\�x���!=\��4#z�5��b%';�'Ǵ���:���#@�9{ŻC�q�p��lzk���d�����Ǎ���P�ݧʾ:�܋C{.!Ĩ�g��/���8�|nS��u�*� е�;2��X�+���	g>u��49Y�*ž ?l5��e.>��t�3H�쫅�_����m��E���M�S�7{asQ��&ߍ�{͛���.+y
墸���׻��)����=V@�kӉ���ׇ� �}�� f'�7�ҵ?:|G�4��U��?���\A�)�����;����u�.��V�{}DFZ;�*ҋ����w{Y�P#���>���9��5�%�;�(ܷؐ��A����cQ�t�M�?ia� ��Kf��ݰg�ٹ}���S��-p��)��t�������ϳ��X��;���k�E~Ї�1�'�N�e��J�?����v�y�}��Ld>�����h�V뉺��pq����|i�Ap�f����Ɋ[�������jL@�vx�6�t0��m<���yi�־H�Q���7�($�Q����NqT"�l��HW���� ��3������|��ļ��B�2��R������_�X�����y���(�j`Oɼu�D�6ᧁU�����פ"�� L��X�B}�R�x՟ZD�nF�Υ���y�i?~1�Ke�n�� IR�]�&5����7`Ϗ��2�����^�^��X]��>���gR�@��.���:��J�� 8=-GVE�^n�L�']��4��T'|
�?����*�	pf��ҧ��~��(�ݏ3����+��=��gjbsL�o���ǔH���Tzu�V9��XIL��a��*|��D��[�9��m�_<N�cyk"����.�3���zw�d�7�d��s#�Z�J��i�`E8H,a�c�*|���h����?5>��-���@l��yp����f�~���d�vM�F��P���xK��luM�{9yyViii�����3�&��չ���Dl����ڹ&|��=cI/����j�
��'|~O�gn��6��,�Wa=�֢P���㕋Y8�H���}����fJ���b�m�?�Q�Ҙ�����?s�u�?���Q�¡P��[�8����`�I��nI�������֔ %Z��T����������t���ks���<��lh���ˋ��.�8B���z��Ƙ��w�����V'����F�]��(��1%�̺��S����,�o���������7yҼW0[|_�������G)�,7_j~���N�)��&<"b����ŭ����)$��#b�Eі����o�pО�7o
�h�!|�*#ث{�^��xXg6*@�_	�_,�2��p>
�j��҇r����hK��#�󌠬��R$���
���dJ�&~�5�~\�6pB�xu�')�os�@���Q�3f��a4k=k��g��}��=�5k�a�Lr^�<�G5`Ệ�_�8'�lW.�&�+LYP#(//���NrPbX��L���\��v#XL�1��CU�t���2�$:>����u��so��0�#:J+�Z�)���f�v�	�U�Q(���f��پi�Ol-����:����.���~����n����=���4Ow^C�����8P]�a��^��[^��6�ΘzW^�յ4e>+{�釄ͦ08ǒ���&�Q�F �p�H-9�UWg�f7؍�纠��6���)��lzb��+�"C�-�Ո�CO��.#�zH����y�����$HS��982C��TE�z~��$�%�C�e�Cʢ7��ق�?��tDy��>j� �l�j龢^,G��{tx�o�{m�s�()KvVz�	|n�#�@><N
j���V�c�׼�<=N�er|}}����l��R��7G�g߿��{�=���������B]��>ޛRZn�ꄽ����ɦfA�vN�(��/��1�ii�y��yBI~Sv�˔��Y#v��fk�xi�rqmq�u�9/�#?���Kv�f�|��3)oҋYG��i�<�����oF�����٩�P^N�Uϭ�w��ę���졔n)�3��J��q�$ڍ�[ݛb>U`1���C�T!p,2X8nC�S@UG�:���d�n�����_C�6zN�[5�)�S�-]���#�L�`R���x���~$�������M��%og�6�ۍ#�r�R�?fpXuuu��hqU�l?�7�����,��5��7<�w�c�kf���Q���<�Ѽ��_�M���0d�/Pg]S_��H!��&���#ؽ���>xLfx��X�U'�zW3E�O�}�����Rm��
߁u?��������]�a�GD`��\w�&o�&W�&��o���p&X���#�!E�~uڶ7�롼���>)K������"y��G���*.l'}mB���������a%������87S�;��F��Gy*)���0)����9��7d�rI(FY�DP��3v6}����!��\�?���L/Yo�M\�
��p��O�
�N=6}�^z4�KKy���\��Ƒst&F�V]�;""����TL�����%a%)�¥[kki	�{�aq��8	�=�,���H9�߽��� �u٠�*{Jo)°! �]{���#@�v����	<�@�s�*(�od�CtA�\?���������Fy��sUՑ����@�ViIpvn��lGR��&2�� d��	AgB*JTN�i�S2<<�ǔ��KQa`��J�J�PD�A��%�m�/jiIx��-�ۼ}�G!]^NΈ¦{� ��^N��D�a��<n^|d���RW#�&]W@Mz�����w����F���vy�y�=��2��Mʏ�<�qk����\B�D��-_+�9D����DAsCV������UC�To�eX��R	��y70���Vu!��g�����۫ et1�����Á���@$�37���6�O�Shy
:��
�N|��W�vCV-D���R��t��vf&ZF�XIiV�������:?�$,�����dO>s�^�ܼK��G="<�c<�Qذ�������W��|-�vv�$�׉��Y�2���X�i��	!����{�m�kx����@zq<ye��)�b��(wg�O�&W�Z����>nv��#~7~b�ؒ�^F����;�{��0Û}���݃���~�^^^^`v:�C�p��<R�������E0Uy�jj�1�zd�Ei�Ztϙ��c${qZ#Ō\p�kz�����Ҝ�}b1����Bʵ��2�)��3�3*�E����������1��vY�2T ��M[d�^��~�����6)P4g$|?�^M����6��X�}�䱨4A`Is��\I��ϲt�4pU��5
<����1@�J\��8�⋄۲Έs�ۍ��N`!W��I+����t�#N�T�$�]Ҷ����=*����1��J[M�E�D� k����ҫ=���E����� ҁ������O��5T��
������MAx�H�s@_���͛�
��ԗyIs9�������m�s�k7��ͬ��r��J�9f91�Y%i)sH��	�[C]�L��� m���[�jy�#YF�|"=�W0X�u���z}��}mч�OY��I2�\�����"�Ifp��P�͎��������0)i%��eA�ǡ|=��Ip*����4��?��p��{oZ�q]��x3vX�סFΩ�SRƟK
^T�x���Р��R�Ē�>Է�o�aI�t��&7yIw���'o:h�B�W������������j�\�۔V-�rwp��o/�&�i�5�JAeef�k*Q?����iao�9�d��W�&�d�����m��d�&��2J�����۷�պJ����V�H��������� �x46�[%n�L��RU����\��a����L�� �PFr6����wUP����ѹ�����?:w
,�*���߷~	��KG_�]�'.2g׋��-%���,`��03��逄uqQbi�3Z5_4��G��y�
��g2�d����#�ы�Ǻ�=����!,9� hj����0�:,�=��f��2@���8k�s<�ܮ�0ނ�rkk���Ѣ��c[�P~����G{y��_.�N��������$��v,LV+�����FQ`��q�";���(�!.���;�|�C�lemK=��;;���d��<�]�2>�����_YXX�e�x���h_ld�[��������K�f@I
yI/
�5\�O P;w! �e�Ka�cxj����i���lҬ�p���0�p8\���Z��=��.�eغ&�o�>1 ,<<�+�Zҕ���1�ض���%s�����P9DpM�E�&u�3����PC!r���%/Ǿ�6`��8f¿�ͦ �+@�H�� ii�eO��v�I���ب6�{�s> �I�����Z�y�Hr���jcAɅ��2&Zu;xT�Oj��A���^5>g����`R�ֹGK�uu�@����F��s`C^� �%�VU{���򤏥����MnI?=�<'V���6�3���Gq�RfQ��U��Ǜ�W0�H��顰�0`��Qc�w�Vb���u�[t1���ȶ{3δ��J~�=���t�)
�jqZ�8*.���r?�-��F^^�Ƅ�GL��D�XS�#�>c�x���NN����Q�^�U�[�����3��h�g/�g��c��"��~䦽2�t�&���"@s�Fq?��L�Bs�.�)�ޯ�W@K/R�����P�(��a�\&3&�B��x�BN�O!3�S��$��$g�g��/Nkik���Z:�bL��g%��Z�﯊l��h�XF��R��f��w`�ųYLI���|㛪3�փ�Kva���R�)|MSKn��w�,Y3����c��Մ<�EXY��K�-<��ħi)��@,��Ot���r1�71eп""XN&�y����o:t0	����z��:��t ��ny9��6����?��]A�aSy=�؋W��2�>�垀Z�NMV�[U���LP�!�miqGg��Հl;Z ?�֮.--��b+++s���;o^!��P��1�
r��~v@Jgz��H��8���a������|<E�O�v���k����*���8썰���;)����/����UU	��Z�����r�3�$������-��d�k��J��G�$a�G���*u��/݁Tx�,~G�S���/ڦ�n��җ���O:]��c��(��,��>�奼�y�ɾ���*h �$�Y�e7I@�u��j#9:-BBB>���,�:"-J�
���e��is�Z�O���]�^[6�rsA��\��&�_�'�,��s���O���ԥ7
�><�M�c ��|2@��A��VP?��|�55�@ q<P���q��2��'#9���B;
(sW��I��P���t@h����s%����aP��2OvxPc�vmwװ[C*�I>�/;!�?�;���Y-��xx6qEaS$����54XQ<�,)@�feyk^�AT54$��=(:�K�+ �$#k�Ϋ��mdl�������i�" �j�4��������/�s�ߐ;�V��N��5O� ϯ00�����y�`Ag��0.߽��܃� /�i���77��l�~Ɋ�����~.�-����@�p�����3�����! �T}�f��~��^��]�!l.C����,�wK�Q�������!�lf���W~<Y��d@0�u��@�U�p��=<3�6 ?Z��.K� \�?7���g���)�����|?T�W�y,t{�$mi~#rUvF\˷���#�=��(#C���3���D��QYH�I?`S���P��誙M�,H%phf�ثcD?jR{Y�����6@�ϴ[�F�m7������G�o j��*0R�SSr�BM����Gt���~~4�>N�GIH�%^�0���m@$�� J�P!	�rKKB^�f }222�����ʥi��`F�)~߀et��} �=f���lj�Xw��C)��ko:��*����tM+�{�z��	����{U�;~�0�:ϓ&hhX�|sG��[��]j��&#L��q2%��f~?v��n�^nW��k�6�2��Ky�f��}b�~���3����5Y9#fzw�5@s����g�}!�y[��C>��в=fi�jj*
��ǿe��|��彿G3��(�&ć�*�.�E� ���o��k���G�>������S)��`+%�J����8��F#:��f�Kyϖ�4ϖƱyv�@t�&��������:4�ݶ,c������V��d�8�7�I�PZ���n?H�Ibxg�`��<罓���f��k�[6Af��f�a>H�����7��B>�{*w����Y*sC��dH����J�qSj@�qk��gE;=�1�,�ТV�($�¶K��Lxi>)Jc¤���w)�;�S�0!�֚���oY��}?��V��=�݋<(�`��+U��A6
�MG�ab�U���4����xJ5�d��4��3W��~����E����N��X��������\Z��
Cɝ;?l��>��^w J�,���:��孕y:���aBO�l� h�4d1��G���Pϭ4����tj^�+�W�Ɲ��,8.(���#����ʢ,�'�r���n/O�h�4��Ǻ���F!1�b�ė�g�_.�BD���?�	@JG��}3�#67��3���C�uo LhqPV�BNN�����hi�����H��
����*����kg�Q����6�֛���Yr��(�钣>,?�:!50�ڐ�4�1�ES���<ξs���{�VvSÖ=dp(�:�:������ӝ�8ˬ�!})ː�7��h��ԫSԓGr���c�-�I�����o�~Zҧ��֫��@=���C�X��fxh��<N���  ��#[xm� IGԒ�(3/b�� q���5���Jh�|���2d ��f�(�}���S��'Y��Ӌe��}��=As��w���Xw
#��/�Qcccp(�� P _6{D%�Q��Yba�&���X�O�3H������{��H��7J�Ez�
S�vC�r�5�ح�{P(,h1A��G�d���ϡ���	�؊��N5�ޣb*�\
��D����X�NW�oӈS��)OdT(�|ρe�ّϦ�غp�v���e@>Y���� *�fˀ%>`Q��#B�G���03-,,�?ⷧ��]$�6gط��ny���l�Ps)�S��E�8��Qm�@�E�>��oM
=f�d.�������3aXG�	�֮}
࿹��͢��G&ES�����ɓ���mX�!�ʉҰբrgM*0��Q��8!{ďf	����o�	h˰X���M�+��{�K�U����E~�F&�v,H�m�����e7o:��=��z���8�{0"�%�r>Mc�X�9�Z���:AKS���<9���YC�)K��۷�\��<�?�HE/t��M�t6�rU�^/9E���铿��J�E��b���> ��,kk�e�2K����q�.b2c�
���ҏ(	�x�Y����xY��|���:���t�
O��� $� ڙ��?<H��{�A���+�ol|�#l,K��q��(�M55�!��X��+�g��Dg&��|�����tz����~�;b"I��7o�s�������I��#�֌:�
H>Es�>��i�) �ȴ!�u9_J&[�S� ja�p���NlqB�jVנ2[�D90��b�F�e����n��yf��y�_q @5yʰ���\�G��Vn���ex��y�IZZZE��:��̯�����3�Zɴ�8�Eշ�|�W��$ ��yl�D���� 7{&�X��J���/�}��Ԭ�w�y�|�g��G_{oe{�;���b��g	#�:F��+�Y:��h�	�P3�Uw����H�I�Ll�$g'�NU�z=�4Ap�$�pxbȨ�J��V����ɓG�(�!��{>�Ds�!���YiG�a����o� �{ࢬs�Ds%',�n���W[D���)�(�_a��t��9|ԅ�f��{�E�$E.�<e����5'�g�f�O܊ᭋMs�=�Q&s��ƽ��)���u'C������7�)�?r���C.�Գ�b�gͯ���xg�؛��I���W�8��kW�y��ޚgsm��c+�K�]����ߺ�k�_����3�fF������Z���M�"�����j��>M1���n7�L/�^��5!4��	UZ�1R�_g��eETN����?�ҾM���|^˖���ՆU�z��Q�Y��U�*�]KS��b�ɫk�-��eP̂���y{n#Y�q̈́un�=���̯�v�����`�e�0�`�V଩}�ڶ2m��wʤ�k{�r�p�[\��s��N��S��-H�*Ƞ�5Ӌ%���׳>b�L} D�F�E�!N���38��?Z}���e�8?��~r�gfDs�Ϟ���Q�δك�K����K2��&ά��k;|U1K�����V�G��#�+����p��'o�ǂ��Ӻe$�G����n����xOB��X�
m����mB�c==�\gn=���?,��5��8~�u�1&�����$��$��#��6�u�6JL�^T�cg=q=k߲�$�V��KH���>�����Qٳ��r$�<����vq�����*iA�q�V��m��{,����l[d,��Z�q�h���na�#@�#޲_��Fs��O�Z�����<3%[�����2u͏2���w����6&�~��8e¯�0��~�z)�D���oM,Moi��M[]���W[�6|T{�̋vXs�m-������;�֛�����-Z׬BW�]z\|��2-1�=-��~?�,|d��E�݊���5�iS�`�e�exU ��~v�����xO|x���F���F�ZQ�l�7ُ���L��\3���Gs��Pٳ�Nt�;lP���6�
!�kx/����e���aC���G�e��~C��5%Y�O9�W5�"����Ƒ��ä��n�r�n��cͼD�x�qrw��y�F��[qqqzL6�0���l��+X���j�G1�Z�M�	��yX�����l�ph5Y�� �%D�P+!�Z+���5��@�b[Sa{^C����:��=�û��m�H�</��yգ�h�P'%+��i��G���-oUe�T����?���E[���V �+b=�%�`5}᦭ ��V���V���]J!�3���U�����(�4o��eJj�k�~CCHƷNfYD姢� ���C�)�3���;h���!Є��)��|?���Q�f�d[ۜ
w�XaV�q�zd���.�@��,x��8+�
��E�G|��M�m��1	pC V�*�XO*������5).�G@^!�~47�00�ֻ1��R^���e*���F��i`��g�)��z�D:n�=�d��ràL+�h��e�	��%ߖ�Z���|��vͷ��ֽR����Z�c��C[�hn~��pF��)S�I�u/����!�$E�pQE;0��"R������i�-���)'g�+s�?u(�'F2%.��W��H�5�	C��"N�> u1.�,���pc�Tj$��'���4�ܛ�5�{����:|��e|�����$�N���l��)���
�G<~���3��ɳ/"_�gɔ/H$Wm]ʻ��N0��ch��W`>�I@�VI�s�eU�{c����b�>�O�?���9>�b�T�fH h97G*;�G2QO�z�]nU����$`�{k�T~���	w�*i�&�YvXS.�|��`+�,\jz�'`{��F�?RHgTm
S2$�(U�M��6G4������ !����C�<�A�q��!����k�f��,�E��m�� K ��:pYb_�e@�E���H$Y�ٳ�0ؑJ�5V�0`��8�3j����[A��`��ݰh.X���j9�c�ݤhġ�.�nQ�*�3*V��s�<�:`�����J�۽�H�<$m���.﨡UlJ��,�M��c;�w�aqD��w��?��2�n:å��Wz��/�$5w�|
UUmL�X�y���ȴK��u�8�>l��8j�����D����UAo�zo��{;�bn�sr.�&3s��h�cʃ�h���-vBȉ�%.����>Xt��3Hh�W��h;w�2����57�KKƸ(u���C.�Dp�D������\ ���.�:������mUW��e{W��86�Ͳ�ƣu���Ç\�8pIop�=Մyb�]@�/���a=+���g���c��9�m�:�.f?a%O&~�J�1_�A����0#%�<_Q�TD�`cv�����?�y��~;^~�3� f?{)��=$W/�گy�6��4�D�H��յ)�/��EΟ���P-�>`ViE��?�ѳJlz�E)�����d��5I��Qu%I���Ӄ��y��7D�'2]�����Y��$θ�v�t{5�:5]�q��8A���W7��W?-�:����,7��cr�w�	F8����^`U*v�=���6��&�lN����I�7�~|=�Co��b�=ɢ$���X�Cj�m
b�<p358D*�loq�)�0������{V���Bw����2���Ϸq8��?9p,�U�1W/��^�\W��,����ph�^(�mՇ�B�� �,�������j;d3��3|��`7�- Y
��_ң�nF�"�y6z�o�����\��̞��a�/m����x)�*�lZZ&�1�]/RYc����JM�1�_H *�
�����p�V��!�w[,�$��7�6f���}\�$��nm܏M���� 'Ty�w��z��PRU�c��\�1��_TE�9ݕ�]�*��"t{�wV��I1Ͼ��s��x��!q"ab�l,�����y�y�:�)�MGX �d=���9���GL4Ͷ0Nf�)	� �F��8��\�$D��ǜ��|Sڞ��/BVW��}����К4������1��BA`K�/��.����񉯎�P?���JYv��qY���m�  �.ِc��)&��.�9`�a�w@8�Q �455�l�e�{�8ɛl�G�=�ѷb�c}��UH�C�,/{�����%v�g���	ӵ����Z��R��#�Ϸ�08������$�Ve	�!ч� �V��Z���g{�7���eSkTTT��A�G�0�4���晫�E�^��Kp���1!G�h6
I~��%��h�7ڿ�y-�"�	w��+�"�δS~c�hQ�
�U��N�h�[m~�}�>Y<�T2q]`�5�w��<ߗ�"�
Ɉ�	�	i�K��)2/wQu72r,�u6�ؑ����{?��1�޽�K)��y�o2��'�^��jn|���4H G��w��ق@��=��[Vv`�벇 �?=R|���,�P����2��E������s��P���C��D7�%�v^�1'��	a�$�F��rz]�hŅ@!ۃy��� ����{Ҁ'�`Dyﲝ����e��@~U��Mw�� �P�����j��{a83�|�ѻ�?70�.]�Q���_����'[��V��XZ����[	��t�ӏ�_��ǹ���)�f/c��y~ȅ�D�IG+�E��W�*��(+a�q""R6���\������)'��"��u���� k�����mm�J[�Bk��Vq1E�Xe([V�8^�Be(B���"RK-2#������D�����$����_W������y����8�<�g�Dݬ�p��L$�`Y<i��͹�3�e��ĺ�-uJ���<aV=���0���M��t&��V�c�w����mS�-���k��<�=���^@���WWR��\o�V�ٍr�6�R���ե���\[���6��!m!��ORZ�s4�C�o�o㒙��זe�nx|FBBB�����P�D�Ċ���|e���[F�IS0!Y�����z;r+0g�~=w���q���������P_�����
D0�X�J���ӠJIBJ"3���e#�Jj��Y�N������o���Nq-�QN"���A�?�&,��C�@����v����ɿ���#��M�b�����W�G�Z�����R�-5^�|��gC��:��X�ՙ{	�&�S9�zmɵT�2��p��}��J���:�\}���ŵ�:::�ݲ�տ���,�����8��	c[�>�{E��)�À�M>RC*5Jx�}v'��``��Z�#��j������A}�A�$�S��\4�l0��p�C���64D��fgg���CN���8�訹�[)`Ƥ��GF�\��p���"i4Cہ�؋�g<H���+��S�i �����M� ���d�C�_'B (h +:��hT�.�	8�ch�!��F^2�*LiW�!t�:?������T%�) 3�Q�C�K�B�p�?�b晝PXB�~�l֊��-|���i��03�\�s0�>��X�8����
�un�unc�H�������u���A��������Om6�Ѕُ�����\b!��>d��jF3c����M��=�L���$���"1�$��r��Z(��TN+�L�+�h-GȵO�������.g�8L���4�%��s�廂�k���-�vSB�8�Ȫ̐k���!������@Y��D8�d�r�`�y�������g���� ��%;i��Ƚ[0�J�끈	1�MTO�o(�Y�O��!q4���'8J�5�H%�7��F����)8d�� 2[�´h� T��Ӈݒ���Y`�lha������VF���0�z��t�Z����n4�����{3����K4�U`)�c��Y#�^j���/��}�Ơ��{�w�w,H�F{�,���a���c!���>���Q��GG�������Pi�.�|/&"t���k(����1:��۪�'�_����(��A��\>Og�4�"�8��ԟ7�'z��؂$��\4"R+\�����hT���"�p��|�;�q�G��X���KkGIk���i�$*�	j�n�W�� ��B�
���ә�	U�����W�l<�"�;d�)�a����Γ��m�ܱ�o�W�cAr*j�k����lnn6.�Q�nf�_��r�߿N������:8L^,��»��Hmx�
��>� �-�0>=�\��;���F5~�v[��nml0=%� 3���3��L��j���]m0O��u*r�#�c����i�����k;�q�� �Ǳ��yi��6<������0;Z��*�9���M=y�����e�i���-@l��Z��`�����D��N��_7ʷ��֤͚��tٱ�����J�k?���o4*P�}�'���]"��H���`ۓ)(��*#7����dca��b�"�>в�(7�Z��l4�����gw��>��qq3�I��v&C���0O�N�+����U����k-[�Z�5�rRg�ʣ�%��Nx�ਙ��kc�b��h=,%��69<6��;'>��ȼ���䲀���P;!�(�� ���T�l� AcŵF��77?�ܻ6���dh]����0M`ֆ���F�[�����öN����n?�\�X��c�6? O�ҙz�£�-�4����<�4�־^Z���A��n�1Vޞ�H��{��Զc|[��t�#�1�[}�z,z���	��z���|l��|�֏��wi�n@-L��<i�>1V�Y� [p��*&�Y]�>����"�/�l�r��q�섄�ڱ�m�sC���|p,+L]�W�h�P�k��h��P�C�����y7��~w4�Re}R�O;��4Q.�S�5bO�{0���*߇��k�L��0�n|��T�DSV����3kIz"����]��'����JP�#m֦��#?��>�J�g]8�8��S坤��,;�	�6�MP�ãO��E��� �2tD�~�HBp���j]m-�� 9�r�Z|���o�,�A;���&A�,fvVQ�L��8�g�a�z�t�t~��@;���Tp���Q���+n]!h�%�joEW��v^�k΂�@�;:9���74�2H�f��~��n�Q5��Dm�����|tUpp�� �Y��U��~��zL�c�� [���Z'yFʒB�~�]>hv&~]X�����7�*����}��Bs	�5�eg��Be���پ�V#y���j���ۇ*	�g���c�r�ǽ9�ǔ,vG@ȂA�wQ2�)���\������PϜ�N8s�Y3���0����������BD��j��D~>����3N�R��u����fײX�q�D���[����N?�D^\�=B�D�ƕe���oE�|���]qtZ+�h�րB�����G��v&�1$8l]5wFy�[�����Ed��T�r��u?y�_�>�����^3���l��ܰ.P�	����j�-� )���)�t��ъRP�=[��N6=C6u�`@�a��ċ��{S�r�\w?�E�	A����X�L�d�؊����<��T����&�H��!�*U��b��0z��|�z�~� k��u<�Mg/iޖSa%�-bs�B���Ձ�d2�3Y��S	`����,���F�:)�Τ�Yw�*Z6%�z,�_�"�ePX.X�H:�����p��4��@C����G}䗀q�(I�N6S��RY*<��>�������Z%K��l ��,0�ԯ��+5~(�V9ಕ�þG�ӽ}}��_�Ǔ�P���V�Mqw��Mbz�� �����O�+��u��N�b�2���x��Č�N��:;��Y5˴Q{�͐�D�$�t"~:�yQ�Q�ה۟_��j:Q�o"0���1���q�a111�બ���k���?�WYk����k1"?�(<���RBy�	�6� �r����N�wӎ�_����_����v���~A�3��(�g����=Lب�wb51���8������	x��<GM��?%�Ǌ�e��A%��,]5��7x����gѝ�&�����(�P*����@��=2����s�z���X�__��ŶHC^?����}�Z 0�ߓ�$%�-	̑�j��h o��:mc��=Lu0pj���cs�������y��~hb���?m��$G�^��`��:���T�_
|����ܶN�	R��t�Gle�B�
�QR{{x�p�LGF�B�sk::~�D{(BZ�O��4��zS�����T�\CK;�
sS��;P��-��Ix@B,E�X<����%$�f�񙗝ᔏ�wb�CP_M.R5�M+M�_���L����!�9�ܞ��~��>����\�%���ч1�D��0�$�_�M���l��zb�r@���;��7�=x�ժ�������|,���mPܚv����P��=����ĵD
��=�_α�E}SS�57غ� ��SAr8��P|3�G�b߼���aG$��?��RR��\���:�@�K��|<OC`3�"|��d�������!\���m4Т��t����C(����g`G�U�fR��0?�F�I��ml�B����5M���}�������"�hKe�^��dk�oGw-[8�
�>����ɕ�_���N(�ƻQ�>�Z�@�37,
�9�������?Cs��zEm����k�L<ܬ�n+�ut��5;4�
�4:��
�"�5!Ԃ柕������*����2�J�>��2y�����f�u���P?_ˬ�����vX��Uu�<����D8∐��� /�+�7g*~�����iT����/���)�6�x���իi�q!-�[h`R�]�6����9s��S��zKk�t�J�N����L�����
(�<�Q���/B\��h�_#y�a�����V����e趽{�Z'���&U�0r�Z�?�^�0�;�*��I�J�Ty�������"u�3�JP�<���E�|�Ǳu~K�З��D6%��κ��>���PU1qV����&��2z�y:l-q-������L$׵�Ŀ��ՒhS7�\577�)ײ�'s�0������c��fh�0������Q�W,�@�M��q�ϝ��I/�m� G!|���H,4��D���$����QPo��4:wD��������y��	��$�Q���X]��H�4��/����3�a5���!�OR��2�Yo���iႈ��*�r��p�`w�m�+n��������7?�cD�:��~�G��o�A�}~T
^C8��w1F�=-!j���7l
�K���V��H��G�C*�:��W�/B9��J�}�Y��-2RWv�R�
�żj��|��%@���N��~��	�C��7�7����7�bWd�O���i������U����"�7��=�W�~?E
��{�02��Yak�/{���<K�У��A��5w���P��qd�[�+ݑֆD�,"�9�,��N1���Ԥ@��1�zĶ ���.��Erq}k'?�x�8�_��d�{�M��m�C���o KN�W���կ�|�i&;��u��)�2I_�	��;2���J4�!�/�Pƫ�����hȳ�q����e���A#�:�xT��p����d���y��@�W(�*�"�/k����h�>��?Dʨ��bJ�T*�0R�y�c�K��E,�J�p7�l��6/�*�-��C}u�U>��N�W��Zg$��rB��)����)}&�{��Q'�ޖd���H���tt������|J'�����^il��}�Fjם�����J�0�U�־�=��Z�Y]M�m@�9�dbu�u�9xZ]U�A�)�A���!?�/�{�[*G^���J�Kk�l�)�	����\�9ad����%���̖_9�KdC��&&\�{?��Z�_O�0ݜ��8��Q�6���ֿ.g��m�UY�zaJ�'��
�V���̬�0,K�����E��-��K;�m���1[%ȅەv��O��!�H(�ђ(��o�b��BY1�r�Z�]m��մ��_p�X�[C�2S�{�Z�s�C�R����Dn~,�8,u���?�:�4�	��b�2j5��|��:�mu�"/������隣8?B���h�����BvE��x"gl�{<��/��Xݝ�+���������E�B`�Gd��սW4��H�_�^�$�Drww'��ǵ��y�
!���
�9u�Si�N�>�͌��%T�`۲�R��k�����|��#o+�(T1w������y�L;-8k��𺃶~���Ed�p��ѽQ�=7���L����Sc���	���~&':�q%��]�w��g��e�Q������0䵛U�W �T����a�K�h���`qY�I�=Uџ�o�<
-"�yf�ͮ�B����B+
�<�{#u�uA��F�a:.)����D^�[�B(�mV��|~D{4uMO�%�g�ǭT��T����\zyo��N�ߪ������!�x=�B���-��0���'�ۦ�5���'JVM���`�p�v_�Hl����hhh0�%���m t�(n!�XE�Y�^�zKQ�M���S�._�~�,z�AdT���&1�az~d��ߝV^���������X�@C;�7��\,�����3<Q��Oi�ܶ> �;�.x��a�~9ڄD?��z>�U{�t��in���ߦ7�����V��f�.�8�yv�Y&�dQT{Z����C�Z]�8q-��X!7�E�!�
�4��N�5�����D���5Jb��\i��'6zN�K�6�;5=��\�޼l]�����޾x�,wT>/�ez3s�as���ZZz�����Sn����\��c5���r���0�Z�*�NT�h*.T*��Hԃ��w��[�e��Z�%Q��hB��ʠ���������-(^Ն/��Rs���~�D���-��a�&�~8�*��[��#Ճ���ric��k��3������ @�B�̺:�2�H6Y�`(���T3$Y���'����/��*�hn7}o0���_T���چ1�m��(�#OI�슀�-��Չ�6��X��j�n3���C��꤃ϫ7�]��)�%�n7���I8ʂ*i?Tˢ-J��[eZ�Nx�5Fs��Lq��o�?��ZX�Amp�NbeY$�1Z6�:���i	ZD�A�?�ꭗ�����wsf��@���`ӛ�*�#@��23�y�]ї��o�4�2������aAs8z�7w���}p�u���H���0�������=�k��T�k���c�O��|m�o�t`��V��-��}� �������:���&t�p�B�AP>�����tz��h #�(�- �������EŠ��?��g�p��~�c������ s9pâ�����i��.�b��d���J��l�NH`Q kb�l(�TƲн����L*�����x���;���ܚѶ��OBH�)SpI��U�tUx�Ҕ��b\%�фE�&E�ɬY�@`���n���D������]6�a�����sb�h�Ƒ�p��g������?Nx�}��A� }%d+���a���u��e���.�������V��i�7�4�vw:%�����S4w���|��P�rpۊ��:��q�rS2���k�<<Z�`�,x��m�?0�18Ȇ��[��"D3�4��
�}N��ɎU��o8�c�pb�C����S0�FifGI_FS�e����⊔�,_C���q�N��^�[:�3^p�`���r8�OJ^:[���&�h�Q��gL-��k�����U�7	�.���E2h��hx�e{{�'�^e(�3A#Q�3������I��7�`:�;��+�>C|F&�u��w��8|K��=�.�����`���OCz��[�~��d�	m*3��^ȷ_�B���=�\Ж#�"�"o�}h�)��4&��m�;�T�����˷�:)�=�_G�������/����M�cW\��3+��w��b
e	�FK#u�M�)�9�k_�9��
P�Y���~~Y5��4��&LQ�+��vxF�4�+ʢ��p��=Bg�e�UL;PwmG0���u��	_�zg% �-P}�>,0��W�����K�=�R����ή*NK��<ڼ�����?��P�=Y��Z��gC�kX��]*I���ù`U�͟ ggg��������!�r'RO��^�
;��hC�7&è��LQD�-L�0.��?��k�$�U:�E}�/��Y/��nͩ�T���y���+�ڦ- �@��Hg����>�z���~�]�>P u:��,~�����ջ_�����gm������~"2�Ѷ�݆=��A��:o��d	����
Ԅx:x��~� H���'BV% ���ߒU�Zy��*M�z���=LII/P��C�������n����8���	aOum���S����g���l���,N
3����R=���M��c:8��,�q���g���������~<v>�p_aq�#�������bu��Z�ܳv���"O�@�u�X����CE�I��Nr���X����2�%Z�������O�\��N�C�꠽��+��Ș��|ְ��F�!��*���fK�W�=>�J&3���m�݉O�T�����8�=��h��~�딻1J �wo9���A3�f��t��'�����w����Q��;�r{�q�'�---@~���̲A3M�P�>wݣ�K�=D"$pj�A{�������^ ��mN���
߳�
0O�?�c�ַ���.��7�,Gf���J���%U��K<�8xk�k���"e��,/�xIx�+h��V@��L�Tf�s5��*�z4toj���J�ފRoވ��ΘNd����:�'�x\� �E�!�)`i@����_��UQF�7�l��� �����~�H�9�F�V]���W�0���k\g�i`;���w�[ZXS-�
u��v�O�c�O��7Ό�����V�K7������뷵��:��#۸Z�����XAT<jݑ~�&�&P܃�-��7ދECg�e������t��7��h�ó�Ī鰫T�I>*ǝiQH >�c���7L���_~ROl�(AsTZ۔�suh|B&�2 ���4k��d��؋��X��xs��*��@���-��>�5Qo˲С/>�2��o 6�Ǡ[�
w.��'O^�`O03�����>�ѭ.5�\�^�}�*��S���6�GRW,��"�}�5�C�`K�d{�Z�t�W����ք(����nƉJY�Eo�,�9~�R@���ɪp���b�ql(o�^a�ߌ��L���u��'�޻��
S��U��]�}� ���9��7m�띕�MrdI�c|l��Z���н���_��FM �|Վha/��r3�XDrUֹ6վ{��Q�eq�� �9LU��#�:4}ы���>w������s�1_?1T�y��W�V�Z�z�h��Жv q���c���ʬ{�Do�����*��zX��Ր�Bj�;=E�UV�a@Kn�4UHh��N�k�.�/���C�LgF`��hD����DC�/��b�#p�J���OZ��?�Lx�1)}�}���U߫���]�u���`���m��C��{3��@;e��v��05�<1��4��o3.&%�Y�!��N|�A=!�=�}��z��w֯�����9�2���wU%@��j��|~�iϿ9j���H�:�/s�`����� �XR�.�[����l�D�� �Y ��SC���9��SAؚP%L�)�hn����C���h�f�է�Y���')�p��^����B���\��W,ڲbnr�$zKJJ^rrQ�4�tל|��K�P����i�O֔�o���Mi�p8��S?��O��?��u�#���R��-4d#��~�-���۰i���,T����gY����$�I��yݓ��;�+p�R�����Xnx�?��
w���iIiNk���sգ�83�yf�g��6^K��2*"�Fbl'�N�����d!��-�7m�_?(��	T�l��:1����}{��y��D]*@Ď�S�m�d$y襒�	#���B�h@h->�y���G:Eg�=���1.es�"�[�������T�Z�԰�w��P�k�_wM��ȣ@�^��j���eM��D��
�+d���JU�0�p������"Ǭ�-$�|�Sl�U�'\P}����FP���Y|�Y�qYx)��͚*ܖ:50}�+)�O�g��0�5A��PZ�}]s�]�>u�i"���4O�@�<�)Y�������t*���l(Iќ���RbՊE���"��"�L"mI�e�����C���Ӻ��:@D����^'i��TIkµ���_-�$ďߖ����v����e�Dr��ݯ�}r�ӰS��?���T�rCjM���J���	��E_���e>�IudrY��{����^�,�Z����o����M�}թ���u]�����6ہxx]m�ۣ/#��t��=�ww��m +����&��+Xq��;�J�gU_ڪîqu��q+���I���G-�6�JԎ$Z�ΞO\ Dm�Td�D���6O/��nHU��e+���[[�D7���x�տ�;uj�-9^<D+�Ke:V�������ĸ���I��o�L���#1������9o7��9���_���!C�R�����.�3�>���_7,V�����M�VAݜ�c0�'���c?v�Wz1J{��m�(%�� �x�u���ؑj���i����mN�Ϧ��V�ҥ��i,BD}�{*C/�h��j$�!��+2�\�P<٥��sL����f��;�o�☿�鈏�_�`�bK���9���w�Od*���eo�}��N�u<���A( m)}[}v�b���Ũ���\��'o�}=e��^�
�w� .S�<���=����x�͆g��8���F�7�:>���;S�5"@k��tJ��������H�뚜4���Jb��>���r�4CD��R����[6�[��'#Gn��'E�>3���L��x��%[*A&c>G&���C�n��t���qg��t����=�i����'5��eKn�Z�H���d{M�p8��������=��T�xw�af�I.˸k�ϫ�߾"���x??(���B�>�'c�2��G1���7,|b#��B���'\֠;��ʻS/��J��2}e�j��(�l�t$�{�� Ó5�H	��~��sǙ\Y���t{G����=�w�՜RXh6ο��,���q;?_��e� 9�)ҕ���	p�Ӭ5����&�&��_�J*���S]x`��le�q�����LHB�K�Y�l��ZU�_���e����Ճ6����>�� ���2��,���Q��ir^�-y]�NW7���`%((��VCY��Ϳ�t��QU<G����&�i��BQHԳ�Jf���:�5E�`;L�tM�/�C�W�$Iox���V)F�����V��l�����d⌓�#�7`F�o	�g¬9QKp��_����a��JT��Awڸ���@,�&u����A������s�mԤ*�V��9�_�wrj�U�[O=�aFzP7��;/	�:���������dX�U�3� }�Fຓ2�.�Y9z���᾵��n"��4�Z'� ��hh�m��}Ι���0p:���mē�2�I�ϾlH�Bh�kj+�ٮ?�2~��"6��َQ���.
�?�4t����q,��r����V.?�9���(�ij�����ACÑ�}c�]���瘧Sj=�j+�R�UA�kc��T�`����@bh�4�X�~�=�t'�u��N��y�-�͋�(y�!�b���M4"Q[CF�u|�������c��vG�h�w�<��c��qIj^k:���KD��w@f�L6�A�������6����-$�퓉�����얆����U�΃]�k7�����Ō�R�"W��<�"��l+�8�C?C^�	i��9�M��f�6�_b������/3q#BVt��hǧ��4�BqN��dӃ��Ov�9�{t�EF�E���}�y.�R%�ʶ�Ҭ���7͊�tו�5E�7~������l�|�ŭ/�<����aP����M�|Ҍ,/g|�o}M�֛%T���c5qʱ�sK�Nӹ�h��ࡎ~n��m�^Ʀ�i��9	�qf_#�x�o��ZZ�0��\_�{X��|3��@���_&�~4��u� *�a��~��!�#��X=��QQ��u왽7��X��ֺO�+����P��������Qs���^�j>{݂��.a0����{}�6�} �ĮC�4ٔM!��rccc�z���I��W)�iYhg�Q\�x|+SUU�P1���ӓ��`8��?$$$<��z+Z����H��JuAX��}x*��|�m'Ȥb�Vʡ����+�٬H/EZ���s��6F`�b�_2�m. r�y�a��L��v4��i��L�e����+W��'l=��o߾5k�+��8�����li���e{��4��2@�Y/g"C��E��7�í�$�Y�J�����ԦUJ������v��\�'�Qs��=P��}�@�g��J�&�)�R�/��������˗/M;��/_�����䟿j��K7X�bŊ�Tf��/U��
��d7������"լ� �k���F��Y���FD��b�ʱTs1x_R��9z���#xQ�֑�qT�1$1b'�9z�<_*yN�κc'�ܕ�����|�dg5��51�BHM�>{��OG�s6����s�	���a�Z�;{�7c�t�e��������8�$�MY&`�|=EqW�����~�����oh05LŜ�������
�,��s~Xx�V�}у��	໑Ɍ�!�Iԓ%w$d�qus���~��=�� %T:��6HiX�'�.o�#�~ͭ�U�qEc��������ں�T�J����j�M{ ~��^����[(��4'�����]���ǍN�/H��(��gȦ�'�;��.��('llk�=�3�W2��~I�!�)eY��[b��>��C��TZ�iE������|�����o*�ne���)�ɦ������A.��P�]}} �s�]�3��|F�l�����|�j��h4�.����k���.�ʹV���B�l�/�qʊ��)]���1�[���ЕaH��妫�4Z�,�_Ƕ�����D�|]�J�rvs�^��Q��)�X�ŋs{�Tj���9��{*��� ��$x���n����l��1~s���A=N�.�xw]��r5����ԨL�w��7��q|�f��)�ԀK,vuCÒ�y�Ǖ;������֤�
�^�z�-�Mq�![�Ls"��*�=��:?���>a�]m�Wr?��� IM1p�A�X �PyWm�ҕ;�f�W^��X}������۶C��ʊW��X^j'�t��q��t�%^QI���.�l�p�p������������J��]^5ң's����S��05q���A}�&�������yte?�CK�$�)��-���<���'�KyxZٴ����v@�oC���QHs���5�!��h����q�H��u�p�e�Mg���2\��;��yxx�r�>��?��s	󾯟n�ݛ
G����������m�X�[d%-����GbD���Qu�v6�\N;� ��a���
+
��t�t×V�p�;0`�^GDb�V�:H��ȣ���]S�����\�p��6�ޱ"�d6Ir?XE/��g�;)��/�����v:���7�"���-�T }�'�$}~���.>�����]<=��Θ��9'�m�%B��b����|?(��~��B,󫱡�����jbv�W�T	��G��5(���Fǥ��;�y�Q���]���Ԯ�{��ج�2� A����J"x��3�u��'ƦD���,�{���uТ�c��cn~�x��Y�i�u􏠧PSiYhT�|Q�?pS�����x��T���?����>c��u@��;�bA���v�,�1G�a$��w� M7G���'���,9�t����	�6s��]��p�c�%3�ԧ�l�7��;m�n�ן�+=q�8S�b�W��U$�W�(`�~S܃}������c�E�`�hd����������pG�t8[i&n�`8��*��U��ɑ�,�;��d�#����K%� ��Q� �%i`���u��gn���'���s��~�����׀e�~���}��D�iNj����)�E��k�͛�:jR.��~>�V�d�Q�$�TtѶU�}�̚��"[̶����9�O8�W����e��{����Hm܊�ʵۥ@r 瘂"��*�F�r������2䇹��a��E'�d�
�f�mQ-G�wƴ;�>2#Ƴ���w\�3��a�bT�3�j3&���7<\�z��\	),��+J�%�����	�RU���s@��3��E|�g�w/W���z�.���)Q��ė%�/��9[ŶA:n[;z��]-蕸8;�p{�}��v�O��W���E- x��-\���!�sl�òD��/.MEz ���ٷo�Ϩ�Ե�s)����#4���a��k���77��� �P�|���q�\���!��A�Pd����Z�٨�?:���bB�<$L�0�C�T�L�.��=t�c����̽���»��膭[̲Ԁb�������a�
���[�m;����
|���k���7���^���W�,ƖE�i۶nM�9�@ >�ROw��rf��Yq���Iv	KmG��n�7�������m�>p	���Y(x���UdA��ߐ���Âi5�E������M7 �<�$��:4�{��~ �G�Z�>>�B�&�ݗ�X��P���4�mͣ`�E�D��h�"f����{o���}�������].&����Y�'��j~�ُ�Q���ywx�J���!7����Nw+�d]�����B&DYEܲY^�kϭ�<UgY�H�+t����9x�.@܆�	�g��o�9y��]#�֜��������K�>����;P�u���"���9d�Z�ӬG:�z���1ZA�B���"�{g;X_so�{�'�~�^��K�_�P}��C��^���2O���EY�Y2p|Vxp_+����\���{s�x�|+;;;N�l�=(O$)�%&�Yn2P���+��T�!��V���bP�-3i�O?���9�!�O��š�T�ࣲ�t�۰m�j���qG(~�Nu���xF����S���P���<g�r��oN�c�m��ץ�(�v�ӌ����M��I9�z�l��4�Fo�TԷe�7�T��Т��x��K�o}}�E�6K
����A�λ)���<����&��m�sm�2(/zy���������G$�R�/�[�0o��4>���$4�^��ө�Rꌭ��U��������3��ܬ��>�l���"I�w%���y_Y8�F���]]�J��RQW�	Y�!��sn郘I���S�B^]ml좹c�U�(W7�g;]�f�UIS�Q���Y�b��Dq7Q��L�{���e�`;�c�^���|�c2�RXe�K<�)���޽{EV?�Al����B�]�ܶغ:�//�\����r�g����v �}pJ��ą�YM�����A>չ�^X_#�)G
J8�L�3m)���Ke�Y�<���TRx��1.>��j��]/^<y(J�������-Z�=��Uk����6B�O�^���kIIH��E�����a�W&0]F��p��!���q^�����)vm�"m��h��e�F=�b2��]�/��c�E��gV��TF)�(>Y�,c��/��S����wL�X:/ύ��|H�"�u[GP@�+�r�6�!�-�ї��Io�ޭ��=%��k�o|3>yiW�E��|Y>������X$d�|v0�h|�#��ǋ%C!i{��P�lK���j�wB� ,}��m�Ԯ��m�w{�� G���m���ٝ{|����n�����k^!z���O�^�`�U]eS�7�$l���Vo�H�`�iS�1EEE��f��������!��ʿ�.��=��b
e��}��z��uSY�,j����tb�TJ�W7^~������*��w�N����8��~�����D�q�qv�@m����=ԁA}#$�mӗ�j7c��S{[(�(����^��E��u�mv�e#���Q��b�Q�,+k�W/!6���Q�Ԛ��1�.�Sh�����F(3x��k�;�QWڭ�M���kM�Z��n>��䍇��a��Z���a������"��7���Y��>��P\Y�v�h�O�����BI��'�����Yl:0��/<����|Z�rS�kݑ@Q=���������~3<����:�K�K�����-�u2�m�.��[*Z����##�u��a��b��@�1�$�gG���3��{��T5��ʹm�����օ0c�
:�A���XH�z��-`���Ww�m�\��R�d�����:G���n �oGh#\M���
�V�,�F���m5����uhm���A�߿Z�OA��}���if_=���c��*��NĲJ���Z�&+��iH���e��e*�;98,]�SہH�8��<E�H]қ��u�]!�ɓ�G�|5�0v]+f��r���~��-��u���u�ZTԝ�ߜ^�ڠD1� yٛ� �5b5��ME��I���nlj� �x��P�����]槒��3��&���aH��E������px�F���t�F��4�PY~�C]�Zr����:m��GU��d��VO�:�\/�$�픚A�G3-�$I��vW$O��5����L�4F�C����É,�	4@��g('n1���%x,D�1w�"�^=�C�.	������q6sW�������nt��s�
�l��dok�"���A�5�,\V��n�w�L�����yEZ���P���1�����ƃ�{xb�v�*NI�SV��������������8&��-M*ij�����ԩ=�B/)'����EA��d�m�|W��Å�Ȓ������}�z@������F��ȷ�Έ�~MuY���#��G�n*IY�r%�Up�cc�8 iF���VĴ�Me�B(**Z����	~����2�#|����,u�
.����i?�F�O���0��u@&����6Ǉ@�P|F���E6���7�{�o?=�3���xT���=�o{1d�l�GF)�w_u&U�P�E*�n�@��/H{sg�_E2��oI�Hh�B }C	�2�ov���3
_�-&[u�R���s.�����ki��7$A�y�'���CaOȾ�˅n[��@��}�m�Z? �1�]=9h��p���O�ff�?��l;.��L�������9�P���L�&�`���ŋ	��Z���U��7];I�k��Y��t��=���r�p��P(�6��=C��,b˦��k8d�=�k�0� �yxxX�Il���Q�A@7K�mI�Jo��=�z��%�Q��Ą�-x5͛�������
t���0�⺁��f�m����?|y�D�Rѱ��;�t�)nz�A8$�6�����h���
�Ào�Y1-T<�Y�e��򾻬���ܫ�K갋9շ����M����ON�T"�ݜ"hA5#/����1��V�bQ�z���<"[q�-�_M���2I�j�S���W �0]7�:}Y�N:�3�0� ��9ற�5�k�]��?�IӃP�^���<�@��b��gZ���ADۂ��ZO ��M��$��h������Z��ۘ���Ρ!������� =��T�uj��&���#4�߬<��7�9���W|���Ŗ]��2��<C���î�ғYL).�X�tم� �2⾕�9Q�,�&��ūV�.�,j�{�2�	k�G����9��:�KD����:��I<�?}6�ś�7o���KdjNL����Q�ݩ�k��\�B&�����kp��t��m��%c�-�V� 5��ccc/��Ի�Dg��0u����8��A�%벗ATH�	E�-�'�l)�.��I�K�y�~�+O��#��8�J8p��A6T�ȳ�V֭�xDA�`A��pg3�.
"N���`N�[ʫVUU%NK<���z�����b>!��z95�ͭ�~��*>9�Zt���]�5��R��H����=����z#��`��
2$,<��,����N���1˻�w��N���Sk��{*\�w�ء��PP eh��ŷo�.d���g���yO8�S�T)Po�O���U- 'c]����ܞ��.uq�ҵ_\8�������g��!�Y�I�p�4�'�ɤ?o����Ҍ!�v��J:�^��<5U_��O/ߎ�塁 �^�܏5Sʍ��&�r]7�;�U	&O4H�9�0*9��<C-w4�z����xP乹��D/�Ή8�5�������B��j�Y2?0!�穦�{-���Ua���r��\o	kO�o��Pf��%�H&)��A����,�⩬�����e��R<���(�<�Et���|�qZ�x9m�r�6$���n��"D.���ݳX��ǟ�?V����O��`����-�U��"�wMk3�����-y�v ��]������ѣ�t�����O�B��q
g��tݐ�2�:�L�b+�����S:�L)W���Q5x)A�FE�1�V�9�?�Va#Y�nA�_!��/�1
<�e���;4t$$xc��e�2֚Ӥ[����hV�_���q|dd䖋����*=E+�n(��Wc�??g�Z *�d�+roMq�3[Q,x������8���)����q
r����9�KJ�ĺ�/=�s��V�kj�0��//�TTR�b)����2�����(\Ԭ��y�]f���c�������"9�W��]dqS5?'��ao�^mS�c~³y�������޺��&;҆ī�I�N���VX�z�UI�	|�T�() Ru��,
N�{ MŮ��9m��z�ut���n�VN,{[qcqU��\�³�d�w���*�-ySE;vhG})�&@5�w?�vʕ��C�Fy�R���^�u���*�v�!O�}�8g�*�#n1������jy՗��ni>�:nQRi��4,:,;��r�d?��z���7�(��k�j�+X�M*��t���� x�}��¢�:28!S��}�ú9 �l!��6��]�@���N��y�dւ�j��N�����a�*�V�b����Uu}�i��GF�j�3=�`�� �E��s�q
w��}�zː� �ibU�����E6q��[  5V���lB\dcS:������+UUQ�+*��a�X ��++�.�ml)O�C��;7�m�K��Y��Aaw_ےy��a���@@���8n�A5�l��֟_�A^��?gfb��aR��t�M1ڙ�	J�G[2>�>�9������;ېr��.����{S���8�d�7rRA6��k׾��f���U �/^��t���Tn!ԭ��Ϧe��_�_t\~h�3d��4���y�l�m����.mA�e��%�)
Ҽ6�?­{�ĕg��b���� �g6��^��s� Xѡ���Ï���Hq���-�Ÿ)NA}����gth��2��]���m�9/W_lqjF?��6�ZK����0F����M�\��k�D�tQ\|�	#�����~k�KL=Ft��n3)�̫&j�_KL� q5��Y[t3l� �՞F�k�����+}3N�)��m0�������I֬���V��76����(,=o8/P�{����(ƙeL*̋b�7V������r�w�5�!j*"��E'�Q�q�v׸���c���_��8��^����r��/�/y����~�cΉ#�_<�bժ�
%�d���[H�����~Z[~�����ܿl)띌Fw�">P.Dr9Q�?���>�-�;�<i��L�����A(a�;�r��`M�Ԏ�ԩ�@�7_��[M��)h�b��N�-䶜V���#�My�
�����Q���|�����bU�ng��9M��}n4�!��E���M(4�)i�[s��W��hѢ��οm-��s啊�"����9�6{�Ϻ�0��}�|z'4�F3��^��^=㘂��Ą��w]�H�x���I�/4|^W-i�gv�x	|�ј��6�����)��l��Y4�
g�R� �9��ǝ!a�������<�) _�����������ܡ���|c��K�J���,[<>K�����U㹭� 'M����I�#f�����z�Ӣ] 8��)�\���h�����m�=N�᱾��i+�Mq��D	u;�Ѿ�\!!!a.կmG!���y��}���Ɩ��ْ;��.��Z��~6��'�:����u�����R�vP���c0����MT��9f��(�
��ʆ-�&Ϲ[�N5�?��<����n{)�"*����eE%BD�\"C�21�iC�d��=T���$�N�,c�-1�h�2��yu�����ߟߟ���u^�y��<�y��I�d��Y�߻a�bt�����M�:�4{^�.��J���9�������Xs�1��� Q�}��V�����0m9|�䱮h��ẶHЂ4���wIv�\���\O�*iL��ӈӾO�]���9�w� 8A]����������G�4��fD��x�i�/��nS��#��2�pK�|��H9i_�G$�U[&k�W;g)Q���t�� җ\;���G���{5��]��S۬��?��~Y���oYX>RI�D�[��x�<F��USx���\ԕ���e�ӰJ/�d�XmC^?*�~G�����s �ЙB�=_��*�JN����n�jL���~�"���p��l~E>Sk��Uҷ�֌d���!u��[j�w�0.�/�+���N��= PMiҮ^ell\���P7��'��i���$x j�\l1�+#Ds�z*1�-��Z�<�y
�M��G� �C����fc�
(#�D=:� $�i���iZzzS?hnį|��?�_��ç��F��e�����d8�F�~Z;��#�7$e���Β�T@�ɛf��zE�$M3�f���a!ϟR�J�6###��~�q#�鑝�N#���?�>OG�/ݿ��E�o;��V���0���U{��Ĩ5%Rr��P�����nn}<'�p���ˡ�fdb"�~��B��G�j�~�&����Ã�J;�0�������5�ۄ�����Iv2R�����Ӫ2��i����,;���
�#�3����j?о��)�yH��M9�����l<h�(�	_��>����o矰�7�E���R�o�D��O�~���0�bo��3��.��ܪ�[L���P*�yu��X /��c��^&���B��_&�GFGW���u�:�|%��6a�XX>�\����|���!FJ��O;:S?)S�$u�@�y&����yc�t�?�� l��u����B������w�jN����N	�|�~J1�s(�;b��9Ǥ��S���c*�R��E��H1�/�����Ϸ�7)��x܃��s�-����r���z��X��S>ף�t��կkM�}����Gt"�5�������O���2���mC[ˁ���\t6��7P��^)�7'���>��= ��ƣq@�����8�H;�a>�ݾ{*�Q8����Ko�k}��z�$]�КĪ�K{ !��-���;�sI�`ėm�>h|�vN����%M/�Z��"�o�=Nn�t7������0iu^��I�������Հ)��P���܌��}Rzv���]�0�.u2�6[=�~�<F���9�֌0$�J�"O�ۯ�o��p��\/
IAB-k�[q��%�B�Ӱ�"+T���p��>�4��7�:;M��[]�ӯ[�_F��cդ���׼MƦgg���*+�,v��o2~�7<�B!ctfRbb!\�n�0�+�U�K��a�n�*cR�l%��5�:WJG�^��B�o?�d��GWD��:���N��jc��	�gX�Pt�&��|��[S�$]�����!�Dk���9|�碲r	�w�T�xow��Iy�a����������>����_r��~�vQ.���|�#O���s��\��
(>�i���)��e]����	��Ke�<���	�:��"��J,�OѨCt<�;p�ضg'�v���y�{�n��.聺�1Vn3�D
n���>����1�^q���_��[ ���8p_`��
����.`���:�6hF���/�-@�0|��o���O��W-���Hڂѫ.g3~��P3�8�A���]�Ky^ywݢ+wK�Iy v��J��Cؗ@�q���ͱd!���Q�����M�WPЦ��*��z�F���l�8kw|���0U��Ð=o�����o9z>��u4����N9�W7��D�Zk�^ZxPf�wF'�DH�e��;�x4F����KӋZ~;�=���N�=d�d˥eu�ʸ��,�p� �@0|-�,�eOo93���^0�A��.Ve�;\&[8qbgH��n�'o�����6Ji���9���v�?��˗RSSs��p;��H��H��d����ͼ��s�y�����Y��	L��&��,qKӁ~Y�!�3N���,�I�
��$�#�>��0�G��N��-�ͣ�U�����RVv�}AV���䴧ha�ӆ������'�~�+}��/�#q����<��.���U�G���ȊS)� �m`�2�Y'˗`0�} \g��P6�����4�$�&��q�h��h�Q���	M��o�5F߾�|������X��վ��N�8I5n:�o��o
�q��*q�ϛ0*��ν4�G7��������mAS�i�}��zr.�]������1�G77Q�QY/!t��;������e$�S(�Ӟ�����d:���N-U�x��[ɶ�1Z7ݍ���~Rơ_敖bB@YE��;9k���?W����:���Y�!F�0���R
��"�'0ᦉ�D��#��ڗyy�4�"�ݷ�Vɉ�I�ɦc1�z�b����ݛF�^��֡��� �R�	���n�C��F쐐(�8����z���ͺkb9���羇䋺���S�!�G������3eɥkQ+W,�t|}�\��j�L�v�\�T�\��y�?ȋ������,z�5���s<��44�LԇXLMJѱ��/@迤���}�ZL. |V����z�����`ʮm�� �C���^T��;�������@	.C,�_'�0�sj�Rp��\��؇b�Cѵ�#�#����f��-���_NLSg=&���C�*l��YtH��Q�8�����df���P���\�YY���~v��V�����W}��=���nnh��}�&�PV	��m����Y�w�N���P4A�w^"�,�kچ}�e�L�7q=G���r����g�h��_�n�0����NCض�+���e_
���^Ot�b��q��\���:#������PP&�Rj�H�8�?pQt��g�p�����K�1gO�3�*����Xt���+<!w!�[�4T>]�$�p��3g�8]�7�%
�#RC$P4�%�?��9������?TؠM���u8ŢS/U/U�Uݔ�����5��ϝ�55կ������`x�Fj�fN�n��+�ؿ���� �n���ﴲ�j.�ptԳ��3
����7p�*'���q;����0]��<(�GA��W��K���%&y4;�W�>��t�S���d&@Z��ؙ{^c8L��j���n)�њ��9�5�)`����ܰ���/�u�t{�2D�)焆$tGJ>q��������V��0p���5TAm����O6����g����s%T]�sa�d�AzW$6.�����������@�5\(^8M�oA���.<r�tJ	݆Beu�Y�g��|��>0s����'����CCe�GՅ���h.�v�NM�����)�Jg�k�p���}]������	��X�$�E��iT���'XgD����-�ɰ���WQQ�{��$b�^�`6b
Lu-�vW�t�DQ���100��*+��#S���.�ą����Rv�Y����T����{�T����Յ]EI�3Â�t-�
���Yl��q��0`S�ԩ��^�vb0�V^=��:*#������S[m+�E3>J�7��qc5�XhR|I��g���,�r����F�s�lv�����l5���B������xH%�g��xN��B��R��]���D��'��i�o�Ҧ5�|���Gqn���' � P�z$Y�_�qqqy�j��_���P�M�/=���sGr��b��<o7��Y�Ԅl�����TF���\#�D~��I���_�"*�ՖbƓ�w��M����C��~�ʀ��]iM��;:�*+�C���d�s�ٽ�?ȶ�U�Y]����?n�s:
��������6쑌��+A����"s����B�p�:�(6�ݬ��nz<�(�Q��U,�9__N��ZO�$�j�A����5P�f!���,��N6g��K{֬��n�UX p凞���2x����"�����c��C�;�f}����(��xV^d��O� �_����<��k-��"X�DN%�����(_��@�O��*0��,�t�DW^��y���I=,�l�-��}y{tt����fJ�B
�T�@������
�!Eg�5N�/���Q�Ҷ�8cۑ$׿��a8�W���1��I/�՞&7*�����W��	*N�k�#�ȵ�"h��k��k��D��N ǃ
�1��[���Տ$MgQ(��
U\�S$�.�����e�����o�D��?Q�m���^Tg�e��b�LT__d�kv��VA*��8�׸�ĝ���y
�ыa��?]�C�"�qM�%x�S�Z!PSRR�8?�憃�Y9�c���{��&�1�7���j�g�W�3m|�[P��ȉ#1R-ǒ��Q픦�&�����~c�Y����LizP�"�^YUtV��]^3�^b�M3�!�����#��+�;��e���
㒨�����9�O���l�bN�GG��/��lL��P����a#���j�վ�FN�m�rֽ)�i@���y�5�Jg�/:���e;y�JM�I�##~���_�L�4�H�#��`{��'���#<\fr�6�����Bu��	�w֑�}c{.]w�jW\���>z{�
�~III=��U}�N(�$j
���\�����jc����
Y��`G�+�6ZTɝ�Wl}�>9�� DJ�����M�*Vք̓l3����Ti��G����N��9��as��̛��Α��
����P��F7��ћ��t�����\z1 {�����1�,j��H���|�����:V�0��r��$���ϟ� ���~�>(�"����9��싷�vm�����2�~Or���$�S�z)I����%.M��e��Ӄ�{G,:�-� �1��ռ]��%�R�G+�a�hN�c6�w�8+��CW�Ķ��e#k��53�J;�[183kcgU3=�Y��ڭ}�g׉m_��:��a|�ڴPp�iq|�^�6�z�OT:899891�X����k8�u�_[/���#+��ι�ɺF�i�m��$�\��jY�=�������3Ƭ���}�RE\������j_���<����ˆ�3=�Ś�Ì�I*I�|�lu\�������ۉG���נ�P�V�M�Pg~;s#��۷ĩ�����E߃J�%+)���]�|���]�d������������{C��1.���-'-�Lu۾i�E�|���J47�失��m)�7(�zO:}��|f�l�K��u�xPp�I>vQp�,�c^0�m�g�,�> P=���C�\�-��m�k-ʦ��tE�W�q�F4vV66MN_=�;�	����`�dƛ*Wx�A��*)J�%��m+eXd!ͣ��n�N�� i���I�"]�����[�d��]iBUhO~��QV�7�1����O��}����'��H�,�-��g�R��$�NO�q��T;�]�j��#{F'�h��6�S�tE�S���@ݧX�+��FĽR���J J�s��0֦����F��u޺n���pKx��xJҏX�F%�l�%�P&�Qx��ۧP��U�{Y��{��4
5j$RH�l��ϋ�D��<���"bp"���4	?�oo��#���_�s��������8������_Cp���7
ʇ�����V/���i���U>L�!�}]�|�-�I�Pb��[���~z�3(�H�٠������h��F��@���r�n|X9�Y�Q��&}������I���$��Y��ol��0�����ni���'�h<I�-Kc�}��[kW�?#`eG$,��9��7r{�=��p�~Ǐ�忾�r���>��j��9��R�^�j	���������4iII����-�iԱH�BZQ�ً��O�t�-d&�+ʌh�����_Hg��w(�ZdS%Z~kΫ���&�bqk� -�T|���b!ؙ�]�[�sff�R�!�l�r��]Z���S*����G{��N��Ǣ�׉-�X�...����T-"����������1�������k�I��Sݖ����pp�,��-H�XF"'�lXô �N����h'�K��Q�ߍ�?~�����	w�7n�MY�`��<	XR��j�!w1F0��r�*�-[���Z�Q��&
G���3�]c��$�>��FvC�����v��f"��zi�����A��L4N�av.#�|�~���Ç�x��~�
kHѽ�4"�k*Ll�%c0�̑J��/_�(�`��CC�٤Ǌ�{2�����~���3sW��$�D+*8�!`�F�Y�+j}���Ƈ	6F=�����{���\���<��"������}^�o�_ً�3�M�Swm����<A����R��ꪪ2� �p�	y�]���1}#Gxѻ����T��OM	m���{_;�ɤ[!(�-u����7֨�����Hzƥ;��|d\�y�}�X�f���Ѧ$��R>�[� !��Y�Q\�	��a���M��Nx�M�H�4g�7����n�ϰ�a��G'xmp.����)��jKIF��uD���ԓI֓���7�� 8m$���J�KI1�����J��LoRB�I����@..?����PK���q**����&�q�b�VJ����k�.5XvG9gX��Ɩ����
��l��E���@�M��h�����v�(�o z�mV3��Xof]LLL����F�!�g����r&�5�*���� �lWfgW��M}�ǻ��FC�4}Ksww��	<���
�>s����q ��6~A�@�L�X��v��cI��O?�:�������9y�ǰ��q=w|�S�Ǧ�6�B� �y�>.8�tM�̥'�A|���D���|�yG7�e�J��&����ϷK�G�1G]�/�(�F�cU�s�b�nL�������6>�X�o���'#�)�H�mi)��Wl(����6z����;-yJ@Q������G-�R��NS�1�-�g��~�ڥ��O��FIf���{V,�����J��/%��zۥG�ۮ���{����Çw�7�F^�~�֍p�9�3�F�D@z�RO��������~��X�C����ѣcۻ
�'F�2��Uk1�d�/�^Eʖ�C��3zF]wr��c��5������Vj*����`[����7��FEe�@>|Q'��,�����Tk\n��ƽb1@֩i���#��q)�{���_����@�
��5�|�HE����ݜRO����,�x�G���`�$�ʘ7F�3�R���^�ü��֪�����$#�-]Wt�A�)+ C5�^�-&ֆLD*����@�+P՛q�n�w����D����~W94d[�ڢjMu��n86Y���^�]�?]�΄��o=�0�}V�����̷WԐ#}�)yV����s�!b�������"y�-�3v�}�M�D}��V意y���YGDOP>�L��4m�6�R����������+�H�5�Pz�t�J1�W;�ܹ3��\[��S�,q=����V��j�١���=$ z�����I�%���W�����<'�_�Q�V�g��C��,!u.�۾���Z�D+�3��9c\���� ����@,����y/-�����i���ǐp{ݿթ� �١��z"��_Vtmi����h*�����? �r�!Ah�t1 ���%��!������C��HFd #Y����(w�|��|�C1P�[��&U��qJ�SnD�QV���&;'�Qж���-u����(�^NT����|�|�M�|���5,�EΥo��T�J&�m���Zܱ
?��6yZ"ɇ3�6YF���E����K߄���4��B�]�R��<�S�EB�5��lͶi;p�smDR[}���*ɑwʜF��.bv�ʕP��'IY�r�K=zTW��,��r�*���i>���!�Dj��H���i�O܉�g�T�&7ɋ����~`���ihh��5��^�ύ;!�����]����B'���6����,�y��>>��e|��Ύ�������� `x����?C/~��fPntS���>7��zD��4��a��Pǖ(Cڂuq��
�̅ޱS��RpP�9�rqf.}k��o5'���u��:&&\r���0�q�['C��Z9��֕1.��m��u�a�@ �?xy5�m��Qe\�Ɏ��N�)l��0h����PxIq��o��5$����!+Ev�]�'�_�M%�www;1�H/��UWlO�Y�ϩ�H1ғ@]l��e9\�<l^9���ع	��_a\�E|��n=���١?q7��`��/Fv��`іmmKyy꡸�ۈ&W��Z�=��Ӧ��P�&�Cgg�E���B��δs�?���0ZEZj���97"H-Ο�5��ok�5:�>���?�5��mX�H,�����
���8��B�ﰺ�y��xIEE�]�i��ȹl%�3��K# �0�e�"�bݰκ���n�Q;���3� �U�$�S�N=7ю�waΜ��Y�� ����v�曤WB����ݞ��YRT����A+�����?C���E+��z��.��T�PO������3o�jf1�@ڜg�,H���<!��L;���?��|b58����~�R�bȈ[`:�-^�O/��s`����|Y���B%��7=���a*7�T��v�'M���Pm����X�E΂ȁ�H|@w�ŪTl�72c���#/�vb~~MY�ͪ�jk?a�(V2H������.h,�8��d��?�ȋ5xN�t�W���^������'��OϺ2���L��A~yW�'đ}�>~��3��z����d�71��Z\���c����-�C������3.[V���J9��q��!�`���uc�(�]Q��WPṷSD3*h��eڜf<���jq��
E�R����ӑ�~�����Ր��
����v��g˝���Q~ ��u}��lKqZ�Al���xE���-C!ok_���_��
A@5��?���s	n��!F�[h�y�W���`P>,B��L/����9V�6 �s�^��ζ�3�|�f��`d�B�==�[\����IR�~�]�"��g�i��k�
6dZ���~�Pwh�8�&\��>ho�ˉ�(�!���{P3�'�d�D7v��h��F�$7(�������rnvf��@~��UM���ʐvT"�'�t����i����a��w�����C��2�k������ @�~��*r��5���U(���ar���%�]����,����&�$�_Z �u��`�gQ�Z��Ģeϙ�wt���e�m䗒�p��_�Ȫ�t�sqv��>����s�]���L )S �V�(}jɅ���2�]%<-����if�S��l^c4�s-A;��46D�F�F5�����3A=%�V��b 0>:!Ё�_2߿;�h~��=�1���.W1g�׮|~���Bގt�Q��[�~�N��7�fG��LorJ����<y��Z�V�H#y��&��p8�9S��F�X�q�-~�4���Y;������;�	5v&�g��*���N�������e��'}Wo�h)��x8|�:��ğ�jqO$�N;_���1�CU:����Q$|�����9�� ��=T�¨�J������6F-��4na�Xr�U����lSP5(��.�!8��A���k�~�G%%Gć�Cn��?��mh��ͭJ�A� �2H�c��ƶ�����^^xY��t�׾Z�?��?�����0@��C�ߚHZ�5l +��Bw2����()��<�#g?vc���犔�k����|?�s��+���'ι�}I%	���u�ۺd�?��!�ʣs7�9�R|Y*�-�ٱ79�.FEë�7������xL^���KQ%�.k
s��+f��vD�[$���q�Ug��΄}�4��j�[�b�G�D���5�����`-����T���/͂�w��[e-�E��yg,�N���w�4�� i}[���j+��w� �2���.r��PN��"�"Q��gs��痾\���8��i�IzK~9�c���W��?�"�9�g���#O�55�=���=����-����Ha �$ :��G�]2���?� c2Kю����L:me��@���$v�^�yuռԟݭ
Il���F�:�f^��As����]��㪐�f9/'�WV��"�w<k��lB5	8�}g��%��i[cg�y���b�#=��B@���Y���8�ؕ�O^޽.��>����)Qp���ha2s��ݾ�����!�/��C���Q�m@��&7��Z0���0�#�&m!�?�H:�)�!�^z2�0�e�����ש4�������7�[?�^o��}�¿�K�'�M�y�q�}ci�OY�v���
���x:(P� ��e�G>�
TL2/�%��Ӿ��E$߿�����[��L��Cf��	�,{s�����o�,ܺ�v�P�
��h�}��@!AY��v+����ȑs,UoT����S����c�`���ՒԴ�����@������閿@JZ���]����ӄi��8����ȫ�݁��Yd<�oRZ�J��_�>��G	�q�\@���n�e2��̿�?+'�*j��j�d���$�C�7ڮ�/���u�K[��<����5u,�/_>�و����i�F>�+#]g	�)(ճ?L�O�Z~5A��HA��k�����؎�t���k"3p�h���ge��\��ƹFY|"l����{�79pF��	��?��,�gh6�ni@M��Xi�l��[gju;(��P��Y��eh��܋ �q�"S����a�1Pb��w{Xy�),X�$��.9�ׇ�R\~"����e$��w��3X�yA�K"NU��y�Y
�x��3YU�a�j�*g��xN5��Ν��~�Hb#��"ը��r�"�L/sW��"���~C���?��i��Ov{�鼇�E�	������P{0;3s[�S��u�z-��n.x��j��A���?�V[���Px�^��"��(O�c��EC���
K�����ș�_�% �V� ���}����xrncދ����������|Y��i���i/΍U4f ��@�����UPfN«.b��!��9EC*�f�\I��Dc\���Wuy�q�%B=G��H+�T��V~4*8s	�ѽ=
`��*NN?��K;H��
�<[1�:���h��?q�[~�	Q�dsC�9�Q�'kZ��f.h�T�L�۫�rx�ĺ��D��h�X�5��r�Z&����ļ�`�ҧ��SV�hTH�iI�o�i��;6���]��<���5ʁ
|���J����
��LOYY�ųgkRT�Gcg�M?֤�RN�$*R��n�K>i�(��[ � ���ת��q��{s.�8&�����W;=�U�L<#��#��S�a*P���n�8H5#�B��~�U�7�f��O6.J��,4x��=z��8֔��������vY-��/��Aa���V5��X7o{�겆KY99;�����{W��]u���^縇�g���vR�'V��={�A�m�Ҙ�4����V}��䟕��FZ HO�iw1��C1�QU�k�`Xt�xz��.ϝ&� ���K����������3c�6� �&�*��� }��J���_۽�4p�/ ���&p�����n�@�M�$3nKH<�ӧ��#��c��"����m<��0x*E���Z��ɋ60׿
�������|����c
��Tw>�	ʴ�nn��Z�I^�p#�������4���s�<)lrSC��W d���%��G�h���I�5I��P ϻ ���|=�����o��U�[z�P���҄����A)12@��zג�ݥ�ڳ.��U�#2w��/|��(Ԩ��k����3�������FA1����+�s��𲡡3�F�������8�Hv�^�[���h���;����w��$FH�����ZC#Z�(��:0ڔS�$�ӽ���k�����:��k�;��hlf��u�[T"�j�W�|=���4ע��5K��E����e5;ׯ`��#R��IK���gdB\����d����4��?�&�~��n��Yj	O�I`.��(}4ZM�m�ȼv�?�4�䭉	��.U���Dty&}����;=��V��ju2�A;<�UGc-wh��, {���/R�����+@�~�ǡ�|46�����*�I� DR�T��p�x=B��P��i3�����:�D���~�w�"�Pjg�ͼ㴇����i]�T��&���i��36Z������b�[Zı���hS�='a���1����۬CL��̑�eOU���������ꯍ��ݘ�J�E��A� t����=`oqc�%�:��0/�WZ�Ѻ�E�x���|��]���$��Ny|��RbZ���G0��hB�Ma	��q�̈́4�C-�Wb��%�n�?��r�ͻe���K: 8��O%7K(@_RAAbW4�6�d:\��P���s�,���S)s�%���of�ؾ��=>3&�����E���rl��;a��Y������E��ӟaS�-PC�m�!.6�4�i~z�@�ha��@����ᴜ�+�c,\�P��(�e��ۧ�������
�� �϶�j��N��Ǡk��'���+��V�^��6�=�e϶�V���^V�G��Y���C
~	˦�#\r���S���tQI��u�*��0���	�3�aA��3g���e�����Qg<M#BV���p�k֔���3jl *�.D��Ed����!k�gl"��<|3_�t��^ڑҔ\w��>g�.���V�n�X������#M���{o�"LG=ۂoI��?�@�̛ر�rX3����t@	(o׺EXb_�Uc���B#���[��;�GO���d̵$�_c�R*���(�<�=��U�}��HO�$��Eh���ڤ�E�N��0�#e���ot��}�~����y�W�I_����t��'�+|)�w�7%I.nd#^~�@:�N�����I���֥�ڕ�_l.����V���	�d;/+���r�����*u���-��?���)��j�"�i���'&��&�����޳y+rX�����D��
������<�<��A��3��-��:ǪUl%�S���¬x���g�1�hB�t�7tD��m������dن�M�kW�!�|�><&�Zoq;̆M�����m=���"�~|�4$�;�n��>uk��jn	x!��?e"ǣ��v���W3Ot[�&�<�npQ9,G�?�aGe��ȣ�kYD��z�a�{�����\���I���H�7!w����fy��U�|�������H�k���঑���ԡ�}��x�55�4w��j�AvTk;���pE�#-2���Uc��D�C'%~�����J"�we��dز��-x�t���{B*��e-��CQbn�IjdDOW17b�R�}W�WU݅���h�oGL}����Np|�EGl:��ձ�G�O[:g̶��œK�}V^��@ |l�[� ���`���U���4ՙ���[��ˡ$��F�%P�u(�9;;g�n<����=���ʄl�̾}�۴��w�ލ�_�W���d�1�E~b|�H�MbUډ�M�O����j})�t~L�`���_�$�FU����h����T3}����Q�0�z���������7���R��D��y��@�_�#�k������]��װM�zL[ ��Sz0�SK S嫙���n�}z��l�~�z��}�`���C5~k��z�HXU�Ƶ����֦O ���9*Z��x���U>��}�������U������()��b*�Ǩ���>�U������Z�)~�5'rX!����@����i�O��/P�������T��<e1�0O�(2���� �"B�t������$YK�?+�;��=�DH�bz�^��@E���<;<1��x&V��o l��NM��[��UW�\92=�EE��7��T� Ϧ�j�7Q9���ׯ_�r�����."��t�g�+p�?�C��\�qhi��Z�l)�-s)�"�x�%��rQ�x3������Q89���I�s=DCs�]O���V�˟'޽�m�UT��D������W�=̧�m]t�D�i�"B�5T����T�C���OD��O�v���K�WU�:�"���PJ4f����tdS�3/���?ga��q �/Z/�d�&�g�� !݇�T��+U�{�Ծ�*��7վ�� N���d�>g���7o�
�]�Lv/S�sq�9@P"���*�[4c(��D�'�j�N�"6j]Cug4hu�����@������nl�ڗ������#^V#,a�Bn�h˺��m�aT6�9���_�fQ��c��u�|���P姳�g$G�N�$cI�ӵR���
Ʃ�w}��-5��C�f^&�O�5K�jO�����S�Eօ]w�n�<g�#�;"�NШ�J1k����.	4/�A�X�:š��,�z� ������F.��Tx��F���]��:�"��rQ� �V)���G�_��Rm�J�����Q}�.D��qu4�O-Cmc��E��xMCɪ?���,�#~�������\Y���ׁ���G��d��7�=L���]�-�I���0A'V�}SP��6�\�z�\�&
g�r����_�9�����t��<���M`���v���s�%��Dʷ'g�̞�V��a�im�n�2̀��_8�X?��y�`l�p�NsIwy�jp+�E x0���t���e�
x�G����K{H-&�#yF^���������K�>2�RN�w�K:N�ŋ4v�~y~���Y�����A�y��+;�Rɷ��}��0@�cF���g�B��^�37j�f�
�ь3m߻kfK�C�VV��3���Ӵa6i� Gz+���_FWN�?%9>k�aB�� �� &��r�#��ќd����D-����V�L���c�a��R_NL�j�EDD�W Ȩ}���s�'�غ{���Ǩ�b;>�f��G�dZr&�$�������m��vҶ��;lj��p�X3iJ�}%){2�
�0�μq�'xm|W^��O�!��6���v�O�gg3B��3H���aaj+�}Fk�n�/�b��j��iA\���= ۾�QLt��m&xW��ѣ���
��h}q�gf�YX����YQ�D>�S ��]I�u�\d�/��*�h�-�r���a�TƟG�-��T��V4�Z~Ja��#���9��cdr0Y��i�тf0��:9i�.y|�M�F��f�[L~`�*0������f��0�[�v�� O� \�Ab���v4���`�Ǿ~Y�Q3s$έ�		gN�!7h����Zow���P���	i����HԽ����'O'>h�Y��4r)h${���c=ۛ�k����CW����>{ b�M��@_���QD�su���kW�s�(Y
��$iDSȄt(���ٙa�v�Nև�<�Yd���������ҀJ�K5î��:��#G$?���R�Y&
m��)�Ǒ�U�gZ{���C���X7������ ޤ?疕h�#PK�q�D_xo$��~h(/��F����54*�	�sĠ�/��uA�JjHЬ��8��$�~�K�)féP���o�d�_x<:��AO�u�iWO�5>�;�V��yy�Ojz�@?[��;�6���@�-	��j[�)�]��	W�O#(���h��M�o ŵvs��`�/���\ 
933<k�BkC�tlk58�E�˪6*8z�[��������T	i�sl�r_C$�j{F]���w�[ڱ�"�����Q���� _;��i\x��JD�ד,>��"���ץh7ۊ�Fr*^%����xI�4;r�x�Yb����v=��W��y�ٱٙ��jPo��ͩ��i䚹��V}[Z*>���A�p/��vM�yeZ����m'~��S�gQz9{O믌q!�EO����`t#���N��Q��N�� �uK������~�=pQ/��K��G�Y*_M�Of��L�|�fL{Q�/��U���r�moE0nx!�A�Ͷ�8CtY�,��Х��%��X��Q\�q�#ׯ��;��6�������ZD��I����b�U�얕�d����(��L;���$$�ep�2��9i�˱[@st��Ң=I'��NE`{��y�g�5k�:�2m֝�˙�e��������H��'�:��ɖ�*I�N�cuaEF\''�q̿x�@�J�9��&�"R�IHj�iCxP�o��A�
��=~�a��\,��%�z�^�0���.�r�M�!IT5���nM�75R	��� �0pb�u�F��������`
u�� �G�tf$d���v�̲����#m�l�-����6�޸�P-$��h��1ɘx�u�[��;���4��?����D˟���D�Ъ�����)����m�y z�"����@�*�2�����ck��wuߺ.�H��>���{�g�L=zt�LY>@�jͷ�|G���F��6y��:��g%Zf�~���Y�[m~���RV�׌!=I��΃�ԯX��?Q��Cj�|)-��1c��|	Py2a
��:��T�CA��	|~o�{5��%����r#:.�����T��L�:��+��=�rIp��I�4���9�_9����NVw���=��@LLoeH�|���g>��/��r<AK�V����c\�1��W��Y�ޘ&�H�&��V�N�m��/�0�w#�	@�\F��ڢ�@?�xL.���>��f���s��H.ܺ��fu����\g��ҵ�,ZH���Y|u�tȔAQ�da����#, ��H­`ϥTmJ?�E��~��d�A��#����7�I��"�$h����B����>��[�J�T\Y��Gs��f��l�3�m��*Y��F���VW��ղ�L�m����߅ΗӍ����E<l��ࡀ�i�Y���}���nKck@�m�5���䆻7ڮ��VFZz{qq��$j�~���ϴ$r��~x#�D��mV�4������$`��MO2FBk�߲!�Yx��Lc�a���Xߘ��v[Gj�%�gH�8<��e�q�?y�7��ƛ�_a��/zrv]���e��[�&����ӟl���M��C��S$����*{�Q3]��sS
���S��x��U=N򞹣3�L(��ݾp�=���l�;�'�T��Lo���}�+������=����wF��� 7�������Ƭ��a�3z��)fɝ}���>�� �'Cg�H�P�$E�~|���s���'.��IǾ`�\*����6�|lI�1Y�N�&�H�^��3(�̧��E�%�I_�����L���nD����W��t�ϓ�����~yY�M�@W?H���������q|�D{�߮�����p*,�ȅ��1���}�m��|tF�P��ɱ�ضA�qn����Y�����@A�\�b�kו�P��jՠc��ԩx�=rGc͈������Z�j�nt��}ɓ���{�����PkyktIGr��iw���!=t#��ro"{��hK�T�M��Z��Z�r���K����!&��k���Y�j�B'
����o�����ㄆ���3Z���C>DK�:y�}}}��[:ˀf^ºǷ�ܩM����ؤ���ˤ�H�K�YՔ6���I�U�:���J49��H4ZAJHb|�6XF���:�F��N9�<�蠟�_�2'�ͦO�9ty�wo��K��l�@t���Q��P�����-V��3�x!�c��� U�S��N�1K���b��[f�R����G���m�Y�����Gጿ2ܚHP?o��J;w:�%I���-�R�N�Ҟ?_e&,<<�p��0�p��0h��X�ܯ��uK}�l9�A��|acm����W������*���J������s�V.�0�.�����ڱ^w]Xy�ڹh��`�2��p�;
���QR�Ղ�~�M�m�:�²��u��/�����Lz>3�LA�J��������Bᝮ�[&>pz� ��{����^��0	�]��$:9��ūM����*�߄����l�hnTB�Gj��W��[Go��KXB�,�_h��|>�4����/���P������bN�݀��(���������3������
W�ߔ�~�Pg�ͨ8;Q{�ť������ɩ?������AF� ��A�x)�o�uLL���<��[�7<���|�#_J�`x��W��.~��q��?�Ƙr_�a���=��6�9Ռ�_݋��>W�`K��5�P��@�%h��:7��X �9�~"�d�-��ƪM��-�s>۩W]ֹu�,<=;�f����S���y:3����9cI|Rpl����V�B�][ ��T�K�h$w�ɮ�+��(�9�#q���NS��ʘ��xu����A�ml#}�z���ɪ:j�M����ipn�i��{��9dm�8�0u�z�������wPv�����?\m>/Ճί*N*���⫝�w!`ѫ��w.���*�CHq��K�ō�AK���̝�Q��KJ@_,Dg�����M"����DH*��?��@x@��6��$��MY�*�rޤ�\��aWW�I������]��x�~�;np�G�^�W�3�O�cC�PFmR�S����'��ҿ~%���
�����/��w9����� k����m�^XEPQ��,�0�d��l!�̰i�UT��f�%�d��"2#�	�%#a���@�O?�����ӧO��}�{�k�{�}3���"߿4�nڛ�ڼ6B��՛=�e�����氶m���*��ϕ�F�Xǜ�Ҟ���5�65������Q���hyi��������������AD�U�ي�3�.�"�n��tGȈo?�����S�N>k�P���lo8j�'l�e����s��W?d{Oᖑäķ<�k>-�C����^��W_���?��n�G��8؝��M1�+��A�w���.������� Y�k�=rl�>w$��1�`�i�T\};ޠ�����c�m�H�$+O� =.)됭���P1	�J�d=�A~�]�j���z��6<wg�W�t���s9n}{��R���z�{���f��iq�9�U�!jd���=pU%��_�zzX��+?�O����n0��
�k����5?M��f2hG:g����QCT��UO5Sy+D�t�Lg�Iu�qX���X��sE���[^���	�b�������/��F��{;��Y�Y�+�pu�2�q�I���z�­����	T���RP%�>W�&Oy�� j�☀XJ������
�^�+���2\cC**4��ʸ71Eme��������ު��w����v>��2+R3K��yo�sh�>�(��>%��J�e۷J��Q2+71ڂ���e������"�wD���i��7�n:�t#q!j�����/ǁ*���/�����Y�����'&=�]=vYJ\kN�¡���"k^��%&�B<��U@ȅ��Ax��;�:��v*��\���~=)5]]��ƶr�PI���Ԃʂ *�ѹ��)��$P^�4�8�V�p�BS�9���A(>{T�4PE������Dg�9.���%�a��A��5r��F�/�Eh��l��։r��W<O�m͵Az�կ?o*�N�<l{��KI0�@%(�]l�uBK0I�tv�t7 ��i���2�>Ƶ%󆡩3#.��ds�1�kL.�R59)����K���	��UO��n�S������I�A"['R)#$u�n���{���2���
g�������y�m}1H#ʄ��\j{����C8dȔ��4�;M�ߙtN�yj(�]1���mn 5��c���*��Ƕh�Z�O���S FQ�%7�I]����#���#a�. g�%~��r�ϓ�CQis�ߢ���M��J��,>s[#e\������h��F$Y76O�l���T#:裕��.���RO��I��Ѿ�-9�Xx��3<*�S�_�i帏���f8�	����ϕ�Ɏ㳾���-�Q	
�B;7�X!�Ikxj�C!�t���S�L��R*�[C��w��'?��v2�Z}G�3��ZKJ�熊�o�G������f�g�288��-1�8�t��]]��C���c���se"u�`H����T�?��Z��_���8j�הi!�j6G��������\�tA]V.��:��̳hVj��ԱP.>����TZ&�*T��?��+((���>f�ľ�b�K�=�N���^��WS�����/B�?02ֻn�
y�!tuA*�<�V�#���G��ݎ(�R'\| �#�4������[�j"��r�)���ڑ�+W�k�	�����z��8����`�l5����Pǂ�mv]]"��un�V�Zv15�7�\A���ua_�r�ښ�2t�5m+:ٳf����~-@��
��OYE�X��%����<��^Ӑ���H���o�^�iB�HG���Z�s���E�5�!2�$�l���HL����&&`��(�1�ݫ?��CU�ta����չ�rB�����v^Ea���$_�ż�Ǒ�+����(�c���3ʱẾ�w�Y�y�{s��<���Mjz8d�Q�	X9{ ϓ�J�v<�.mp���c���|x���~বS�جl\ `�q�I��^$�˕�;Kcw8�E+z��/t�U,X�`k����4��+��>�7�#�f"�2\�qj#�}x�S�2���&���"n�cmo��_��/��$�^�"��WR���}�UY�Xn�c2PQ�'t��J_�.\�+�����c�	��2�Q�$@Z��˴}G���W��7{�7$9�負�`c�ٛ�2���� ���ٗ��S�t�N5�X��|d^���w��@N���?pL�m��u�����8������W�����r���OQ֑mۘ��%�D�;�6FՔ��GξLB]�����_o��#~[��%����kWWSc�N`U�(��~͚͓��#��U��=$N�ޚ��t�ϴ&B�I~e�ʒW!=�ʮ(��
^,���]}3�0�m�~�;��� Q��+��H�ڋO�	�~�SD�aU�樂�WY�P�#�u�r�G�f���F������^�ۺ���9�fЭ�.�ȷ��B��J�СCH��'�3�>�O���^>�o�ɳ�l8����]F���|+��������=3H��|yЩ���^��A�d�
عv߉��6��(�ׄM�nL�� ��(H|�.�_,����.��Y�����}�S�e�oG�e�]%w�nn�}cp�����X*9����n�_����Ss�Hӡ B��Eo&�]�YВm�#�a��?PqY��E�C=�������ns�~(�Yh��@wbW�\Y9�9�:�Y�}�Oo���T�,���(�G���mgg�B�;`��!-���:j�2���+��QGo�ȯ������(��☗�O��ixQ����p�Ko��Ԍ"M�H�ӂ�<1�^���(a�=�[)�G�0^�	Ȃ��ti�>� �u,��LV�kJ� ����ak���{?ݯ�m��7mfdj���S]ʄꄍ-�g��i�0;B�E,���y����t�f�]���l�����/T��?S�W����5��� �E��777W�h�s�tN�g�<���G������4>5f��Ѱ�H�y�t���1L�C�$�=�$b��#�cvHl)�k8�n��U�-���cOͺ�U�.�ƭ%~�8A��;�716ִ�I�Qq�xk{;.�vC�7�LQ����?5����و�S���mXSVv�;�56"�q�I��|�>��J�;�P4��hL/��-��@lH���q[p�����Tf5Z��SA�����],�0u|q~���.�����Zۦ�� �mD�c9*��("XjqN->�w-�����k������W��:����L׷V���=�-�� ?�(�����.z":����F'A�����cee��	�f3!�8�g^1�l��̫2��Ϗ�Hk�W
B��ȥg«J�7r1@��7���󟉋Rpפ���Y��k�xD�.׼�>u*��/���1Ѱ�Y�+]��o�J�G��s�/���uz��3�u���r���!���ǵ�k��K{��r���mP�;�(�]ASo������t�5A�96}�,#y(Y"�V�7�:�0#�����AM��H�x�����<�o�lC{}^��Z�ͲZZZ.H�����:�P��vN�=���H�I��D�
�qx�`�x:;~?���W4�[~` ���}aA=ڱ�]>E���g��������4��~�Rq�t�C�yp�a��?�Oç��V���f>w�g�7u]�Z�~z��ȏ��P<���{���͠)�D�$rŲ�-Sӳ����[�2j�5ǥ�z/zD�'��h/��񔿆���+�M�}[�����!?]��(��F����/^�|�c�?���1��ǃ�� �ܽ�8غ���	)���W��-,���N��hE�\�X���t{j�ۻ��O�/,#�gR�,fr��Σ��4s�1¯ԋ�OS/�*'�ρ~�R	0����Y��@���`~j�O��3�L��@�;���T����S?�@��_����CK|>���B���ǒK���^���Ӧ��N<��ZOK�n\HW�-JJ�R&���v���`�t�>}���OF�n�x�G��m"��\�F7���mY�f�?��M�iҙ��YW����ۗ�������mw)��{��H�2��x���]�&=�5�ѣ��B;7�ƫ�,����uɱ�/�d%pa)��?��	����.�g�����UJ�$
�b��xVZZ:"&�9���qz�%��/_Δ]�M!��}�騜\25�i�lk���������Gz�D*��x��Z)��%T�X��6���>�c].����I�RH�GBh��7��G	c���4�l$�h�w�M=���M֥�7o���	Yo�4w����d__��@r,���d�kd��bWi�Z��(;�X�*�Վa0��ޚ�Z���!h�Bӳ��&ߛ�d���W�0���iR8���v����-v�(N9r1��g/U�.�f�����B��S�M�J�+��{�+��>P�OA
y^��+�M1�V{Wh�Z��۹qh�7�$z)�}qUbd���¾�xNS�x������,��ﱶ����?��M�.�����w�=o����I$�ْ�"/��III��56a�O��г�a�-xrB�.jK�,��)o�0���^#0N��U;�	�jr���{v�-(�ZױrJ$��t�����E��իǟ7�E�,n�u�M�)��i���x�	m#Qr���aͼ��˳�g��s���RL%R�	��k�C�G2�
km}zi&h�9� ��\1?�ڼ�nƪ���'�0M��h�a�'o���x�p�MN����+L]��,����������j��ˢ�5� ��tb���w��m/?�tt�ґ���'Z���B�/Lt�'��a�R��腻���d����/���0�ai  QRr򆹧������VVo�|Q��;��=�>�QKr 4��[��W͊G]L�$87�`/���>�
���[�˧�W��,��Ez��S�&���)�Py2T5�n8D����S,ehnj�ȃ����=O/%�O�o*����[�:�u� ��د��Co� �F���־��I�4����(��^w�#:T����!�yy��^O��s��\�H$��ǭ����ohh�[R��Y�h���8:f�~��k�ȉu3�66�`�ubB�'�/�e��;]x��L��"Ж���W_�
�Rh��W�:�A�\��d#�w[����v�8�D��L�U�RLR������́�U��b�l[s��͛��qU�w�
O���=�H�0-�j(�y�*y�����߯�]�7�Of	���P�Cw�dLV^ŷ[G����ȉ�O���6N��4y�1Q�N�+�r���ɱ�.�'��sCs5N�ݯS�o`--U��&�R��C�Q�����?Fc�g����v�V�Ap�լD�+��a�e��r����Q�����PI�u�E��SO���ݛ���Ѷ�GꙠ�n�=����rI�SFEEe��t��pojk����6��G)/�����,�wN!�i�i�-1��D�p��>����Y��0[�����m��L2�!��c�� �5*::�Ɍ}��?���Ȣդ�j�63��Oڢw޻�*�8KY��h�G�@�����Ez�bM�<��C!_@�7"Mu���5���ݻ;h&uutt*Î�����u�����V�y;5�a�<�H���^j�s����vz�䋂�n	t<��j&bN��a����3���'��F�����>wԍY�}8�L&�I����puk�K���i,N�N��)��Y?�5/m���7gZ4�V��+����Y��Љq*�����Z�K	�-�?��N�[�������Yf��R��ƴ���o��}$ā�[�=�����ѝ009k����Q�=��?	Z�K�S�^����t��6#{_ U��+w�(��XK��h���&�珶����Ex9�QϺ���C=\���Vt#?����C"�!��C�<�8.�s�ojN��&q��K.��F�D87��n��;�YZ�L��%yW����Y�n��h��0O�t[Z�st߰cs```�K�}	���S������
�uww�$^e5�?I-cYZ�B�ײ�"ZP?�zyG��t�]�"}̪���#bZ�|sZ�W�3����Ix�]�<N�qh׀�[����S��FFu���%,���D�\�:1m��Q���6�]{��(���$d��gj&^9���Z�j�A��a��e`�ls��߫;�����	,�,:K�ok�m��x:~�_��8�\�����DoSz�#R�aQ�!���n�3�i��=�vց�w��mV������B��U��A��H�'gw�!��t:���b͌��u�VH�0O�l�au��&�_K��d$$p�Ѕ���z���e�۷oG(��A��O�Z�*�աa69�M�Sxш����A#%���{49��&��p	��`E��*���������7�/A��C�?q�r��sr�)^�5�m��گ��=��W&e���D|��!J��ݮ�ql�>��3�B�0����<����h������ĄG����!H{���I��t(�Hx]�m��"">�	|~���[ʸId��E�GG?|��Qά�lG�B���F�Kan�e���M�g� ;�}��",��$z$���>N��3L�c\�����ܼT���gų}�s��tT��!F�mx�"1??�%�Si��׿u���C/�@��یfL�>�Sh$���8�H���0R�y)�3$W��.�� ����z�����ͺO5�g�T\�8����������.��6��~rn�!]"##�a�݇��;�>EK��:�^=�d	��\��#H�>
�ޥ��w6;��79G��z�'ƕ�"��h�Y�*��쎸��֚3��iB�T�烵�~i~�9)'?��E��F�#�#k~ġY/�Eg�%&�6����ΙgH${��֬=�T���6��0xԙ?z�^�B���3�XSAG�����{Td]wp�&Qp7���k�ж��zM:��^zw��fE98�1�wn�����_p�ȁT�E�`�3XC�� =;�j�N�M�>�1:K3a�m]]]��v��*gn���1Q���xs����@jNnn���k�ڂ�C���"4؂P���7|v��d�Fg\�HU�_��}	��u�U��q�@-�VF�<����tꉸ?�j=�-���s*܌n���56^H��@Fpz��9^=(7/�f`����{׀Q�����e�t0�x�b�m����hg��;�@�V���M4{��n� �j��ex�^ɡ�8>e
z�ς�)��0���Fe��y�[FTh!,~QW�f�[��m�逥���h(��׍5�nV�oVc�?444��.�$�
��ȼ�⚓��z+�/aZ����(+����m�WWW�:�KҠ�ޘ�;�@{v�-T��H�!�*�p�I���xo�l�:;�(aml��H�i�E���S�?��'YE	s܃�zЏw����,p�+z��׬Kö?1k�1 �8T�������?�.�mq��Ilm�y�}S��Ŵ�Dx�L
�f�:o��ă��c��P���!�u�����4	z�����%m��r.���d�MM��Ə�8}���
.��u襡ѫa��+�67�^t��hrOOO��~hk�`NO���u�P�z]|�iH�3�孥��/G�ـL.
�v'��ϱ������,�+�!�@���>VO�m��w�_|b�J9b�
!z$%K�M�C'��F
[�RU�Om���f`m������G����/�E��:��=F���Ԕ����5��7��,m�xil�50�UUU�������ߝ�v����5��h�@���!�t��)u����0!]�mN~DZ��Li�D�%�M� ��pl߶�;���"�;P����@�W$[���� �����λ*�׬�M����w������ݻw�cwl,=�W��;�^�&�l������ �[�"�/���3�¨������u�F��L����!H��L�Բn��n����mAX5������j�t�kNkr\�%s��\����F��\�mMssEM��D29�&g`B��U69����$�H.��j	��W����]�T�9">����w����݉�*���ޅ��n))#�����e+�&5:���uxT���wvu��Du�b�c�SRD�
��>n�&�CLOG���P3����ϋ��)���ʻ����B��3c��h��X����.a	#�FQ܎�T|����K�9���5D60~�YV���h1b;G�ߌ�@-�ȵ���l�R+{6~*'�A���9�X ׶��70�yx|a�+@X���?~��� �e���X��^�#F�zeW�4?��n�K%��}�HAUr��j�_N��3[�/���h��rUj��YR�@4�7ǁ-.)�z0�a7H�J>�݁M�{�C���Ϝ₼�O�,���)�#;98�ZՔ7�����(kf��y�됋�a`$��� g�GFG�'tJ�?�� ����WI琍�ZN��0��>兘{�����a�=��txk�÷uv�̷��Ō\����Q����Vo�œI��̓i�,��:Vw�����B�
EE<�B��
D�|��H�Քݫq�ŏ��;9���ZIA@�_�� '����<�������iI^�(��g�]
b�$.���M�&s��aگ��'%4qn�P���okk����[��S��=70R���#��f�7�M��J���WAF�0Lm��pI��QMTDD6�&Ӳ���5��_�y���Gڢ�MU��5���㛍_�=F~{�&)��� B��MM}�f�%�c;�KJK3��7>>>x����Њ�2L����r��	?�IޕW��*t��� 9�3��s�E������M����N���@�G[z����\$��΋�κ��������͸�-�:�Y���u/����u쏊� =���°�ō��Kb���ܛ�������l�v
�C����.��N��`�ag����TQ�b��f߽y�����k2i������J�C����?����OD��{7}g"*$�[�^U�/bE1��r&a@d|�/�+��ۤ�������V�0�/���r����^����oߞ<p��Ҵn֥P� 2u��^�z�ݚ�R�.�����Ě
*�a����@n�Oo֥ ���p6�<�}|�c�c6����L��E�bk=��듔��xm#[��?��W5>֊�;��R>�� 6�fxE4��E��H���v�.�j��@�����h���e��{�]
�U�4o�����q ���3|���khu)��n��C����<�db(Me��4����H�fyg����&�AOnFo�'�_$M��_�xdy1挳
цY�r��<߹�mj�3��Dkjjr��.R�������Qy�<�?�f��
�����R4��Ljϒ��_�/0�a��3~�w.AO����� E0P��76����n��)�PZ�,�g���1�,{68U�X��q���+]�W�����e��k��2Ll�)�]U�l��G9�R��pY��4[�=���v��?P.U}T�r}VC�-��,�}ҒAG�� 	�f,�����gǔ7��f�����k�~������tp��C��Ǔsd>�@�1�Yݟ�Ÿ�����(=�'�����&,3@P��K��N�p����U�.h\s�� �u��*��k�����%Ju�D�4�I�<q�:���	�60.���BhD�w�D<̹a��JL�^�pH�V{��-K<d���GnA��Ả"��;���G�tQ�������q������s�8�|XCS	ʶ���m�A�^��PE��1ī q���(�H(����xג�j��W�M���S�][ŝ>��۾�iW��\��A�oV��#�!w!T�\��q ����^��ޡ��^1�9��
_��=Q/%�x}����X;��)#Lٕ��K��Nw���?�#�J*���~�|�0�<�9���{��>{#��<|
R��q�Y����|�kzǦ6�_�� )Dc�#������I���_�7�?�(�-G7���?#���MWƱF``av�����F� �����\ɺvLz�=��*#�V*��r��i�	<i#��i��`T}��]=�5M��}4ePhj���~2��(;c3�F0�2ӱ?��A�Bti�dH������tDJԺ�$�"���诜j�a�`���La���,��Cx��r�kI��M%��i����	���B'��l�+`�����8C�����s|y*��IL���G>����0����x�ܹF4ӖZ�3��i��rQ)��b�u�$���Joٕ_vaM&�\P�΋��nׯ_V���BH���k�m-�O�\�a�+)�@J�ă��ۖ-��\3ҵ5�Jb����J-a��H�%��S���Ң+{�?��L���L� ����u�(Ȳ����ؾ̨R�
�1U�TVc�n�ԗ����������{�%�F��T%�cB��&���_|,T�Fu&c~U��ʨ���Kɢ�����mT���$Y=&T\5Hm|���@`�Z�y=��|�����`�C��:k�$�	h糃�ӄ.�f��X�ب�;u2HlE	>(�,,�l�[4���>O{j���tSh���7�eb�ߌ�͍o[#g ���<Py��s9������kL3��w ������c��q�q�)]*����}����I2L��P�P��jѡ�WZ6�Fsb;�)��;~�L|�U��ۦ�9g� ڕ<c�Q�3�q5�4�\�t�S�/ݲ^iyd�Ǒ���޴+��`qYfVs��<|�@Nl-����`�<!H�_�n�)c�J��#�4�K^4����)�v�*����k��M��֚n6�μ����II:�J�+Ј�4B��P��..W����RӤ?���m����Uk�� IڴO�Z�'Y��Q@.����@�0:Y#�����l�S���ݯ<�
2'g{AK�X�|f*��RXRkjy�:��C�d[�o����_�{R�W��Q9ӱ��}�O?K޿}�(ao�I���Q�F��xz�YOW��ڏ��DV�� <l���j�7���>o(pb���݆A��zyAn�dy�=�������������	��~��7��q��������djƃ�SB�4G�.;]��C���9���������׹k�������Z�֧��\����3j-�R�̾���!`?�� ��Ԭ�փ�g���#��KY�%d�^�sм�^&��غK�l��t�VZ��G�ciY;;����[�?I�`\1�򺎇$ëpD�w**����`��!Ю��:Q�����?,%fJ�-Ƿ�k��[�$ja�(i[���p�؝x�g�(�#!z�7�l:�m������Rߘ�?����"���5OmD{a�Q��<r��
�����
��H�FM�SE��z�J$��3����,�܀v<���d��D�4�.�B���b�ĉ��VR��������^�1N��y*:��մ�4Hc��Y)� ��)TX��������SGCS�Ј���3�1p�ҹ)�ݝь�t5H"��-hJOt9]��˷�鄛�<1��NMz��S���o��Ib����ϏXǱ٘��`)�TF��3� ����1�Bʹ#јŞ��N�M3̬a��W��͡}4R��+~��$�m��Rh�$K9�o��8���":jQ����՛�ֆ�q��ic�	m�vu�F�#���$�� �p�t�tt��)��Dʺ����Z�����
���������J#o��z�	��W�Q@��=77�g��O;SX�u��;s���"�/L$�L�sѢ˶J�j��&��0OJ����:��0��[��;�y��{�ʔ���@��p���$	�KJ=���ݾ��[��y�H5�$	'C;	V1� ;&�ҿ;�,�Q]��%c�X��؈��^z1�Ϣ#��j�pn�`)U�̜v.�&}����<���J�W\+ExZms90����i��	`����Aփ��t~�`g��L|�E�4����Bdd����d��%|-���������vrÆ0誎���j���V��B�����O�:�c䈺m:t�}T��x��I��&����SG�rN�y�C�G��2�nI��wT�B!�T��^<���7zi����1:ȩ��򔯑t�p�/�A*�R�I�&&��^�/��v�(���C�n?����>j�ϥC�:� ��5@Rݘ[�a�8�}1Oڢ	�jY�F�X������!������\�K���L������_f��zN�.i-����̼ �Ǚbʙ�h�s�F
k����ˇ��J��}$��L���@"\�U�>1�Q�up�I7�{�u�}��\�M·w3w��ןh%~&���<0Q���c'�Ν#�� 
;#�@\3����ÍT�I�#:���þ�7<$�N�U\���|~$����w��2���}x��ݹ��}�{ɳ}���V�1JA[����jQ�@��C�c8 ZH񘫔�j��l�1n���J�oo��2s�� �|q%N@�͜�	�-!��N-���j-�yd� ��V��- ��k�u�ʶ��+����Q@j��W��O��i�y�R2a���Ul��`��#����6*��siO���������H�<��J�*!���~����v��fS؃� �|��_ĩ%b�vl�ǰEﭸ�Z)~�!�g>�D�J�`��� E�p������ds9�7rb����̘y�s��h�s�0Xu�U�vtA[-�w���:m�k�L�S�0�()+b���؜~ä��	�N���z��r:�n�O��ÛJ���7�g����;�s��ՍD�](*����'K����(
��0�y��U9�b�$Ā�&`�@Q>w�.
`��C�~����i1~�=�"�I3�S!�2<2bRZ��yyFcaF˳��!DeWx�F��<�$�5幑���Ⱥd�4�l��j����Tm��ԢG��W�����;>��h�]HLL�����kum�7�l����$���5G�ZoTd�J���3�U�ǒ�	��ml�6������+(<�ė��������~�1�L噃�V��6����Es/�`r�����jk	u�U�O�*��r֮7|V�/z%zx�;&��!D�����,O����rh�!['��#$�#9��KpĶ|*��E8N%�}�N�p���3GZѱl/�?@�C�r��+�A]z;��kN�B����o���B�zE�
廅5o�sms�揪ᳬZ�/�r[W;^����-o��`�ZuW}�~5/>��jFM�Q�p��S��1����R�h���'_��Mٱ�[��VQt�c	��kǦP�,8�Ef~�C{�UN��F�C,�y��g$q{=H�d��n6��f�b	��u�����E�61�V�ވr�ZL�ёG�+MT������~�A����C4v�	ʰ�c��{�t��6]-�aa�8)9Y�P_c�DN"������.{JKK�}�R3�p�����倀ιi0&�66�ء�c-��#P�$'L�Z��3y������^(�w|uL5=.�tH�%�Qf�t�0�Ęy������z+w#U��q���k�Z�\���b_ޏ���@�Y�鏠�#j��`i�׍�������TBe��{�m�<�<L_�m
돲=R+��KLݻjU��
+"k���?�����t�'0�ٚ��̕Rw���hק���~9��y�ߩ�(x�jOŌ�R�Fs0)ŝ�ͩ���f��/PA��.�4��;P3��`���v����8m"����&�����]1ݶ��Z
	U��n�u	88���M��ѳ�$��H��	HT�~s�lIv�oUAGG���KR��S� �r=��S��d���Vl�H�� 7��1�Y�lkp���	��5}�J�)�ó3��^�.�ğ/��V9��FY���B�a0��@�ݳ\¸�!��׹��6������Og�4�X�P���E^����ի
F{a�D?%ȗ�d��{��}��$Z��!�
ؐ3�n�]����;�C���4ix��ٍw\�� �k� �>�Zi����1 �e��-�8���@����+r٧9�Bzu\]h���Ō�����q��̶�o��H6��\�_��;%��	�m��O��Q�E����V����n��Q잛+�?4��`>B�6�*�X��_��&�"w�W@IYYY5e��26_��� ��..�_C�<�`����Y5w����co�G�m�G��M���-�J̐1�3N/]3���
�;�%3�+��o�07m"j�76K�#�a�;�	/Vӧ/I�0��������]�lm��}�6�0G��.��wBU�dP������}�X|)Ϸ��0+J��3R>>>�j��1�H&�+�������-�9U��7P����Gw�)����{�x`4ǻi�.m����	���O�=�]�چ��8`��c�T{y�2�����Lue��!	���O��.6����DE97�Š�e^7:2R_Q9��ԽVSa���ĉ�S���@�<�~�Æ�� M[04F��hk�b��h&�Yρa���K�M�4�H���҅^�C��V��er�~n�-G�O�����m--{f�u��2��
�ύ���_]u�9T/ZUo=�n��J��!���r��������#�T"G�p���+J�^�GQ�O�H6LMD�.�U%��j�:�����zVK��WS�Y<E���q�,l�ހ��j����+4@ߗ?��Η��i�H=��7�m˅�B��Fּ�$VT9�Ԉ��E=��W ڃ�O��iz6���Y:R�Z�ڃ��[���i�,�^�h��sp �(U����_����قu�J2=��w�_��eI[v�K4!�-�^6<�Z�'��\�������%K"�{��Ka���cu�?.�u���Ů��n{NSe��z6ُ�i/K,)aT��&�F�M	`@�YZ�A�|�̟�K��p��K-<YJ������P��9R�P.��\��5f,�[c�|�T$g�D�
�u,��3<Y>�]�Z}�1vm����@(��]m�V|���^��5���Z�/֗+��A]g�Lf
��&�ԍMM'�W+r��cY�X�A���&&&1�ڻ81L�R�2��(����i-��sѤG��ho6Ȯ�7dW��}�˪PVJ�v�-����r.�� �ҰB�R�$��L��B;7�1[�
N�U�u��폵��n˗�d�*��vڕ]��fX�A �	���X9�|�eI�D�Hv�˲Y��ve���U�'؝��Q��T��&0%%zk3zѸ��,:ޕ��A��΢g���WM�ʀ�N(D7Q��Ҩ����9$Lg�Oz�=�-�Y�}���i��&M����b	"U�[��/b[��D��19P�@->�LÑh�Q������m�~eߙ����=����[N�=�h���S��V��������;�ߘ?(H|�II���ˮ=G�cF�k���,W~�J�:4� �h��B�9��g0��k,ޝo�M+�F�^���Rw����ˆU1�.���DJ�K��[�v�zWkw`��K�F��%�W��� R��O�������������<�<B�/�RJjSS�\��w�:��^M�?��Ρx��L�ֵ���)�$�� �17?��h�͛W��bg�o���VR�r
��mo�_U�l;�b\�VWn�q��ܪ��\Y_�kbR\1��#���A��/���juL��[��m_ծ�)��~L�H/�&'ejj*�l����K� (%ED7�}6u��k?���c>&�}�
tvl��g���O�%+��`�?��F ���wgHy��S��.��8�qQ�R	��C��W�����QS��8�^� ��^7;���A���u��=��%o�����4�g�@Q�Q`r	�������+Y3�Aw�`=���3(���:��W�rC��=�CQ�r�g� uuu��Ґ���@�R$��L��cݴ�Bd|#��W����h�<n$��k�մ>���ӍCSY"D�i���Rո��#-��?�jI�7�f"v�4�l���0[[Gs~O�-��۰�-X�B��epp��:�k�ѭ��ʙh� ��!��@bvGU0��s�4��d�D�Y���eW��wo���r #=1�]n��������6�
�NR����>���IH7�A���kG�!8'6�8;��M�=�_�n�y�T���h(����7������sf���U��_|Յ��n� ���k^#�u�x�[��	� l��8�4�3GhtC�� �d���m��$«%K>�[�TH�����*Ԉ��w���Q;��ZI�uE]�}W[�%Nv����e�n����}��Z�o��FB���&�ǔ��z)��ࣼhR$?���"^e�k%<c����s)�]��WFu�����d��p,eޏS�#X�P���D�FP8�ي�z��czـ���٦�\;��֤��\"�����^Rd�*�E&�G�;��-\�H;���C����A&Zu�	�3�r��'���H���/��>nMt�ީc3�8"�� T3�|N����>���+-��̧�s�Ks����}r���H|��O��|u}�����D ���q�\"��u��P��\��J���F�uxI�+)�T{j�	M���eߘ a�ħv&_k�U�����R���.ک2�H�y�
����
F��¢��!<O����`<�;|t���o,�U��bk���@�($�=(y�_����ID2sȝ2������2�kkNq��w���x�u|ka|V��ߴ�.
�O�
V��`��Fgkl��޽�<�?�J�d3i�C��yt$凱��u���T09H���4�N+���:/���?"����p�����>�V\���@�������ؿ��B����Ht,w&��C��Ӱ�"D�Oh�\�6d#/�N3�4�+�'���$1Cj��OYӝC �N�R�}�N��g�R3K �V��Y�:u�u}^�4�8�K�XB�)�b/�U���3vn�:�'��<�$�����!v�Z�KNW�-_u���hgQ"����.�F���1ÀP ��x�>�rߍ���x��ۙ�8]�7��n%�.�#f�N��u�F�ѱ��oO"z瑞.�k��>h��K��מ���b�˯�(�Co��[﹪H_�S��G�3&�H��8:�����.��{�:P^F���ba�6l@�8>>�ao:��joXʢ;�ω������ԋ�����z�i�,c��:��G"k�� ����U�b}mot�d�7���(�c�&"!���<�z��qĈ��/��索�A��޵)�.�~~fn�999RE�?�P��fU�.���>���9|�:v��r�4�YSss�\�4���hc�*tnd��9{��D
tQ����/�P���os�ꃵQ����ڸ�}ҋ���_�g�-l� ̂�K����{Q����o��T�+�[���,�\��\��w/��"+�#P68����~s��x��,u�����4�^Dc*s-�b.��'ˣ*��c���@�u~�*�]���c��J&�6Z��܏�����L��w�l&����u�tg�D�K�����bݓ����i ��3��m>�uI��pI��]��#ll�Ңϱ}��<�=<-�g�^y������%�������!!S�f(Bj�FFꋆ���Yk�����zl���LL\�$�U�u�N����\W��n������$Y�׮����C��������6z���'�����i���dsP��,% #1�p)����C�4���h��J����Đߦ
$֣�ߕ���#��p$�s/ڕ�޿��c���?J@ߨ��A��D�k><H��nm"����F�C���K��Awn����qE�T���n��)?�aq�Q)���ח����5@��cJ-���������V�͖��^N)�������U��J��eH���#�.��Hm�w0���
�H�-��'�F6FP����=�ϓ��𢏌�x�h���;�����|ϧ;I�q��,���P����=�үn�@����]��>k�X� ��>	)	l��,۸��$N�.��Ѥ�^�O���Z��x,���p|���B����Q�	m����B����2{�������'<|��pH�+��S�L���i�7��ơ�׬KՀ����8??��N*O╬��ʺ���Zѐ��f�=�܍k`��Mdv|��j�E
����H��!BmQ@@oW�BSCE^9o$���vM����.M�BbQ��a, �����6@UË���Au���A%tL_}�Ԃǜ�Bzk��.��w�q��~�ZY=��j`������}���.�x5�k�񨦴�jF��E�X�	�Qޠ#�g�G@Ф0����I��N)���������/�͡���+	����QK��3}�:�:��
c���Sb�� ��'+U��TE�.�
�3[�_K�ЦFa��φ�����oJ��J�������.\.����ɚ'c̗x�0_�[�V#+]+5���o��/�+s��@ЕD��e��	����x���k@�8�#A��&��Ě~�<��G�QQɔ,]�c�]��W{��ٕ�L���d�0���1m��ů�&mˮ��� �_���_S��J�+P��t����Ԃ��ߚ��3�WJ�[?3����Վ))������<�T�6<�y&j*��O��-��'UX,�T_��;�2��p��m�H�dnaa�K�0�5"1Q3���p|���c9c�9_M��#������������ ��j������Ă MAA�ZA�D\Ddi�i�%H�  �E\qi���t�^P�RX�9ς1y��{�����X�s��{�{fΜ��X���E��k�'^�`�')$���c���a]��xG��@��'W������ƿ���-&|Mf_������v�I��G�����D�M� ��E��Q��������|͟��9�R�"�����]��e�q�Ͻ,O�~3Ū����(<���4tu�}MP������R�|��X�1�����.S�����x���Țz�]���� >\=pBc��R�tt�%Q?�;���~m
�T�eH�w��&0%����h��ۉ�F�ԣd��p��{�et(����׌"Ȉ�Qj�����Y��樫�nt�{Њj�DШ0��WMt�~f(�@&����JMq��A"w�T(岹��<(��閺��@k�7q�gi�;99=����E�;e�Z �c�<�N�k��.�ymmт�#߶/��
��!�����I�����֕��MNN�q���>�~���.�s��&*j��u+�@rO����`B֎4�����%P9~�`9_&|�O ��5?�! �dcm}U������]�l�����!�&G��	_C��_�Ūcw�� P$�s�7�e�Ne:r@yUz�v�~T}�a�g77# 2�sc�yl��ᅅ~kkk���5�Xخ$��m\z�mNk��$%-����Ȩ(=��1.����Y�� nF�{4���a,�� ��I����[���� ��^�xI����u�_Z�MΫҰ���Qş޽��q��^��|�3[�ηX�|���Xm�����K�	Rd�Z�������	���-���~�J��#�&mâ���E�Ip[�:2�E�������M3��-ȱ_������.��m���6?�KIII贝��l�nrh���Ocl*.iOY������#�,rDj����D�Fݹ<�~�A�|���GCOSN��Q��gzO�����?�$G����C�'����:0~>����`�%FR�u]�!�%#@\�J����.x겫��c	��{R%
f6>�\IZ¯l��^*7�B�d:�V�@ôDx8�ב5�>ǒ��{�K�ѹ���&������;���6n���-��x����T���M��Ol�;��T�N��r�(i���C�ш�2Q��B�$F8�F׼ij��9���R�j�nQ˲％��H�hTX��|�]4&�ekG1r��nmaq��dv��%��]
�m��l�;�eR	�y&���+aUm2gV�h���"Q���z����~�nO�I��t�"R����Q2ލd���q�ٞwu�Xqq�(�S����b�ڮN.f��a:�yrH�f�x�2�_'D1iQ�B�&?.,,�:cd�,yc���N��\{ �8!��n����<�zR��]�\��qLp����G���MkTNj'�j���ެa��(L���h�Zr�>�p�P�����&ܮ�m@�Е�{�z��RM����ϒ�3�?��.�P�;�Tw�.��}\�&�H/V3���0-�-@L���d��dg$$$x�����������qF�V�V�.<:19%e��6U�.f�����c�����R��OG����0��vn�ֲ�M������Ot|�]~�@�Zb�]Bj���O����^�Nĩ���zIu�J�{���զ=H _y`��=gt3m���Bxe�j�'���������a�S���(#�kX�,19
7�G�b$$$�<p���7��b�z�1�n�P�+Tqȅ疢���`J�����h�m�C�Ŕk�@����tR6�>�^>�1��8�;�`G��a-N�B,��eV��,@"i�̤fb #�SəlNWכI-��ϟ5�.�w9�7lڴIQ1�W&�/:�ܓB,]���g9l=�����W^k�,Y�1;��9��nTAAA� �����hp�X�srWtY�����h����/ s�qt�i"�D0J�E��^��I-��g���dO����N###ަ�N��}�K]�TCA۲���j���og��ReAt��hHܻ���¼|�n��@��&YW;���@����ܫM��@� ��[TE3*�d!��
���������{)�M0ݰ���Σɒ�H�Æ�(H=1.999M,3&:�`aa�5LV��J~�L`��]'�g�Ʒ�zCV���Y%t'�f�+�um3�����-�<����G�uD_n�Cg�7�\RfFia�V~���1���֛ockI(��2R0[��%�X�g{����e,�o�?RrI%6ۮv�k�ֶ��;���q�������iW���ķ�:��y,���x��rUH��,�Vxϭ������o]�f�^u0�7�A7OQ�R�x7��;D9^�3ח�y�D>�j f~:f���Q���O��R*��h3!��qW%�����͉��S�e�(��j(�@�W�p5�6�?zc�3�pЈ��v"^^:F���(���#�*ε�(O����d/�m�D_���H�a���n=D��J��.����<wJh
��mV�c����u�Xr'c����A}ck����o��hߓ�S�pӬ���mU1W���<(`���#�Q��4 ~�n�o,��B<��yQifD��0��(Y���>��e�wj���"��-�����yt[+++���N8dG����v�����.�h�ʨ4x#ο5��Uv%%���^���I_Gr�Q�}����)��,��I璼�-j�����9F111�v��L'尾x�����H̫C˚��T�
�����7��
�*M�q��bI����S0N���U0�4������;Qυ�u󅴞k�^Ҿ�"ɻƓEwAGz>0^V;�i���z����4��{c�v��z`a�f�.��h(^Qg�3��Z�L
�����(��;��7m�~b����Y����b��������&��<��c:��S�� �Y�]��>������t�˸^^
�!4Bg~�n>A�|i�/�z�}�H��ިpǎI<�����`�Q��{DcHHH`)�W1�zz�S+T�fdd�ۯ��@�:�Y��͔Zk{oU�1֥!��L��K�ԡ��_�Q��[놌C��"l3����Uй�R��t(3Co+ơ]+�_����21Zm�R����p���;~�׹�ޚ�����6̍~��+����O!c�-	))���j&w��9γ�b��e.��u:V@D��1Gm�"J��e8'0Z�ͯÏBz��F�>�%�AL������.΁?SC��,��s�^s�h���#��{6�2�P�,���3�vjQ�E]>���PMd.��e�MP����i���N#<>�;ڬ*`w���u��燵C|R\�!�u�E"�_<���EKx � ńX	��B�"U�)?t�<$���i����4�UTRr�I���e w��1W4�vv6���q��>����:��-N��	š��Ɋ�K�����M�j��GX
��/Td\���:�-� 4�סR�'�*m�6��;�����IeS��6��n��|(�=r"�f��T :ɒ?��7��܂k�L2[f�:����]]'"""�[֜52z��.ݾUCu{���U�N��Y/@h�@h��u2N�pɻ�U�A�75�)�4���K�%5E���<�ejj�pu:���~��1�u����W��(�z6ӶI��U�D���T��?�LP�"*���A�nn2��A?1��I���6�r�9��uz%���ϗu�<� $U�M�.�jЍ�y>Ti�1��P������I���.�3��(&�,�&�Z 5����i�A7X�.�B�/a�����IT2�=��w����!׉��槦v�7 �ۿ�ؙ+|��'��`'(��z0p�o�-Zk� ��+y�)�v�Y*�`_�u�!S1JLw�Y��k����yO�x��1󳽨|���v>��u���P8�ri��(� �Z�:���%��F1J>�SQQ!Q�LSyՁ�σ�X>z����e����j��6�� EÜ̹ �JW!� ^{�S�V�<4����1 =����NBDB3W/$\�}��"�O��I�����_6�׶O��F|Qe�E�T����$�e�w���H�V(�g��^�$&[?ZD���6�#��Q���Qg%����o����(s���(&`u�M�Z�v���������BXF	Pg�؈)�:�w"N�N�2Ag��y�<�;yy�~_�em��5}*��Kx�К�A���Ϭ�"�_����M�@��:�ju`�A�)jA%��Pp)x�M�ncR!�v�E�ݚ�p��Cx�p-�q�B�#����� х+|fQ�J`�222/<�e���1�(����@��|��]z�Mb��
e�P_�bf:[p�P�r-�a"5��X��%��Tx���E�@�(�ۜ����5�\�u���]g-i������~ff{};��.���Z��	/D;���? �B�nmd熩*߽^��������^�8Q4���+�;���)Gد���o��q��n�ޔ��#]f���67��1,lK��bo�v���edf�,"�����~�/��Mjݪ�J�C��˷H������4+8��+�wm�jW���z��y�5n�֫��u��ϻHNN��%[X����g�N;��56Gmy	K����'&L4�f��w����,`@sC�s�O����ܞ��޾�9�����zE�Y"/�����dbFܬT�[,�}�B�'�e��aE(Q��75eH�5�6�K�q s>�������� �W���%�s6kx��"b��Z[G2��FVρ=�T\\��ܬ�X���TG 9�eyv�+!���[�}�_��;L�vsu��c�%�-�W>�§4���+���{閳�p�Guuu���%#�p�6�t��淟��!:���u�^�(�����kB�Ov;H���~�k#�7!��Q�^���l�甪��^g�Kn%�:�E{܎"�����k[�v���?���sHLLq�=�k�t(XyXO��ۭw�.��ASB��W��{��<�PCa����oF���-zi��_~����#�O�I$���;/w�*�ц���"�/��ݗqa�L I�}UB฽a�u��/w/�T<�5��>�do�.��R�W"����d=`��@��M=�X�y1�s�x�e���[/n�g޻���sG����/��2Dj3�^72b^���������&�[���/��r�������+_"�_��@��mm��W/�##k����R��)��/ ��[X�+L6�ӳ���d4:{�����մ��| �Q���'of�ŉGai(Tcl3J�z�����Jug�y����^):�[SV~��Q��Y��iwR�CRn��v��j�ú$.X��C�
1�egg����%U��t�śp��)�M1d|ʗ0�^GxS�'�6?�N��If��$���p0NoB�匒��KH��ݿ���~?o�Ɋ>�E`��r��5���#����$Wi�/����
�WOT���b'Ebۣ���"��ٙ33q�ק1���)��O�b���/ڑt����h�_ѓ������'5�F��wQX�e���8��zxgt���J֬��=�Wc�<�o[� �^SS��2ttv��I�K֯��4i߉���,A��R���
%-[��Q���{���Em'%7/n�C�h֋]�D�;|%�X��˫}���Z)(]��
Nx���g�<3qO�*�vZU�6��*fڬ��@�2��Z9�Z���R|"!4w��?�S�	(���XNzk��@�
�tE�ȒK%$:�1.��w�jT�w�[R�",2%��N�m��]�GT�@�F�n餖�Q�5�����hb�ò����ƮW�Y>��]��,s6�3�ai�'RW���x0l�K��- �8C�ń�'�ꉆ.��SRR"`UZO��
�����9�c	�,_9�D+���kP_���M���hF9X���L��� �/�y_u����-�MG
ރ��~c.�z��O�	�7�R"���R�"��}��H+q4���,��
|#�;Yks\g��>P����z�5�#)#W��� {q3��(�
���RL������\�2�2eU?A�Ѐ-�v9�_��x���U������֮]%+%���ׇMD13���>�Z@/�v7���I�,P�&���z�V�N@hRQ�j ��C!��IT�3�r�SA�%$$�
l�]���Ⱥ�����g��6������4KJJ���$Fį���<�LWy�K�{��Z+�U��g�ASb5S���C��5��]\���_$���Ƣ���oW8cg��I;�ځ���q�F"���^��F%�̘%Ւ�@���Fb����la����#h���8�Ի�ǥ��tw��i��V��ۅj.46:��HkίVUSc�\��>ϝe�g�;��V������C�S!�W�36�-/W}��k���ں�𣝍͚��e,1r� U�}��ܭ_�Z3>��/���!�7���f�OJ�@��XKB���ۦ.^Ak�n��*Ea9(��0��@^YzI\��ד�5՝�Ÿ����.�l40-n��D��΄:V�+Zy���J��<���=���%Ѽ��{3>��۲���T�x?��º�͖E�5[�4>���A��(!@�Xߣ͞��ƺ�tȺ+_v��^}�����)M�~s�����������N��A��q&[���q��Q�����z	a��6�#"&��]�3��RR�o�Պ.x��򔕕AP�^��?�oj��a�Nc,�������[D"ꆁ�˕����m||�
���ޝ�kPmVʓ������0uܴGq�θ���u�Xdf���m��!w�af��ե���յ��;�i���؋�rW���J(��~���/ g� �o�F�4�p�%ԕ�Sv�@�ڿ��n �xP@"!�����0��������R�C@�#��~���un�jP���b��B;ŏ;ac� t>��}f�ûjN�����%-J+�4��MiX�5��/^���z��H��5��H�y��9�~���9 ���m������!���2�ňS��w���z�����U@���70)�����;5!�5b�����/ܣ���d�c� ��=�>{���L����ؔf(������ö���۰���j1���0���+��v]t�E7���^tQ�9G���v����`f��&%3�b�'��(���I;gz��%'���;�lG�;2�R%�neiy���A�*;fw�X�i��C���*b*L��s("����w���*o����p4�ˈkD''�n޼yd~�VR]�� �3s�G�d���f�;��w��s~�j�lr�m��R����幣3�!��6|��4�d}�=�!j¦|f=Z��Q���܊�Jzi{��,�0XҤ�=�,��*���&A��@P	8�Sm�樺*��,�!YYv�RY��[�A$$'���ﶼ 9U%��w���j��>�0���̙3�(�w,�<[`W��$������I)��n��F�M<	2�xÑF��yx�}q���/}I~���H���S-Q�c�dz�}��c�xTQ��fq�E�ҚW�O�yxx@�Ƚ��R�$�?u��4���nԌ�Oj}k�J����ؠ�z�{W�#������%S��n�ef璳�D:�OJ����ȞN�h�\3^�u�\�p·UIj�R5��5��8�0U�'~����ŷ���X۽�_Ks�a�y����e���+��6���b������ 	����L:\~;5����q�:��� lh]3�s�%�����\��sL�b�W��-�G�lه+���V���W�aMT�U�eee�~��n�vO @����t�bAl
�;%--va�����`%�Z)f��!efB3�x|��������\�`�xLC��k�F=pލ��yK��}0�M��w�&6_�k�.J3V7�y@O@�.�]����dM��UO3|�[�mL���E�<�11���IaD	��ĉ	gy�)M/���\R����j�֒Vl���rr`(CorIu�� H���^Ywڣ�~��C���Ffн[����1�,z��f>��\�H�kmy�'�}*-��km� �œ��,�ܮ�a����ځy;�#��ݪ���C�#B���<b_*=���P���]~���đ�y4��ť���oc���_�|����D���2�&O+��XND�|�p!�O�x�B���!%�Y,�R|����m۾�[�z/�����Dܩ���!�\H{��5 bw�Fww���y�:��F� @8�F���\�^@�����VO\?5��WTTt{����nPM[ZZ�Ú�3��a����-L�L���F�٥ϟrL�G��iՠ0Ndt4�.+����ƥ(?D���L�����X�'�9�h��>�F��f|�c�K[��pn�U9[�����_{{�(��x�f�	#�]��p�q�(O���(����-�Ġ&,
F8���v&贠�a��I�>U���:]QQA�&?�ۮ����T�%��_r��ذcr-b���Ձ�����m��O��	]0600���f���NpeЃ՗u�n݊���x����)�v+�Zl�������ݏ���V��/�5���M6|���l�/��"ɸ�ש��Qc�����g��D�+�Ū/�񞅀?�@�k���E��*u����˻��J�/[�Soѭ�-B"Xu+����%������ ��2Q�� ӵ"�}nB?5���⒏uS�`����"���D�O�>c� �D��R�%Q��z�0�_u�J�yi`$�a~�m������f�;M�FyP�h�����R�i����<vw��Z���i���r�G�F����.��&�H̿�6�AiS��CQ��:��A��6�}Z�v�"�|�B#!SAA��1��|��~=��#��0�dC@�s��5f�gⲟ�Z����{�#�_췻Vcna1��QS��P�`�ao(@��gς�֋��EG���i@E�P��zjٟ[k���>�x��e�<|�[��B�P�x���ZQθߴ�!��@x��B�R��|s�L��\�t`����:w� R�u��|�O<~v ���w^��Q+�y�^K,�?X��.H�X?���߹}���ᎊ��Iz��_-lH9� ��vb́{%��^\�&<�A��-�lW`k���9���U�ς�EyjtO��ǈ7��� ��h_�iB�kLj���1�������6@���'A���Q������z���3�{_Je�DF�s#�jvR> (�M�"}��)� ���:������R(��*��X��;�)T<a��Dǆ��"�ب&�:zݬ������!��*�	O�{��䊧uO�8&�7U����ڢ)Ǽ�v4|�p��n9�r����ߙ���tI52=�t�#����缙)ͦٛ�-��X�����t�QC���w~��N?� o��sxX(�b_P�_W���2����;�m��� ��|*Sq�ż����7���U(�kg\T�
�o��m+�ۘ�����,�_�F3���<T��Va�Q��6�����0��]zv�cE����t}~�
0�U~��׽�tW�>�=�d��J����U��q�������3�`�O���b�?r"(��|�ԉ�����L�S�G3b[�`�h�d�KFԽ~}�2���eT��A�U�}�����Hœd�h�D���1�I&��!ۺ{�cn��[�t<�7�&��N�s���Ȯ�3�k�CtO��"�@H�6>�)0���4`��(�ł[�]#4��oڄ�b�D�����<s9E
 ��W<�%�T�����<�K*�,��1P��&1�Ɣx��8X>Sm����h �|%�{f�(��,p��w-�XB��'H�,d���QR�7��&c�W�s:�rnf@Gķ�Q�^���_����5��k��
���[wP*�o�GM�%P5���C���M�<�"M�پy�D�5��`P�{��EO$#fz"���L�p���z�������B�}N��x�;��i�<l��v>����1GE��[}�x�֎хm� %���?��׺��C��RLtS�Ⱥ��;w�خ��y�X�+{�ej*���۴�s���ձK0Rh	}�X����һ���w�D�$�6��I1��xg�ndh�*����0�*�y�τ���~�_�{�	���g�'��O���G��H_ﱩhO�KY3���'ǀ��@ �H���}JPޖ�b9�*hH	x�1|Ow_<�@�B�����x(B�������޽�u��Z����I�c�����A��������+��5���m���#��沨��;�f�<Z��g���x�_X�-u'[t�R/�z��y���l�Ak��χ�Q���(�{��	����@�֞���c!��s7U�k0��qʳ�8�Iu �1Yg[�޽�0=�?��n��/�[2Wc��;�f�֕���F�K�v��d���Ok���Xv�M�P��\<����)��@G����d��iŵ|
�L䙬P���NG44�3�=���Ԥ|�3��3�:m��o�~�UBB�es{'�����Ŗ�Nc]@�$ �M����4F%��=�m�M���DA���&_��پ���7��d3�fh�x��]��>��n��]ml��M�"T�����ެ�F�//�(�b��u���L��� ~���J���+�#�r���[JH�����/�i��&x_>P�R�;DK�Z���hhr{���<�%��B�(>��3]#����HMFk��%�����}Un.�1Z=�O��w�lS��4�B7'�O]��d(����-��.���s$�[�@����7�B����1�@	Oi�h$�c��f(å�R��k��>"xr;�dʜ�ԕP�%���R��%n�8�2��H� ���a��];4D�v����HEEe�{
b����j'�V榒"�(-�M�dϿR���kh 2ǯp�jQ�G�z5�������'������$������=��D2O�G'��߿��s�(C)��g3m%A{ݦ>�N��zؐJ��聉��v�B) C">�� ����u�B<���]��,f���:��ŝt���$�X��ϭ�)3&
a�b0T
��쥑�B�bB(�@L�i<3�	��T���@+/�mfR��I?�h,���{���*��-�z�mO��h̛U�d��%/��6r����8�>֋{��q~����5�O�����^�hȕ0�����d.?KXQ��N�H����� ��5��_�ڐ@� ~
����$,�@Ծ��p���-�`t�e��̫��>F�	Q��B[<<�ݩ�*�ljz=���e|�/��K��#��[A���;��K�w0����d/��_�@%�_L6�����:���� #1����T��l>�C��6��^L,�Xt�c����n.��k?���
�!Ћ�\���U�۫��W��|�
��|Ƿ�vW�ܚ�l|�L�hH�Z`�P�SWs��U�6��)3�d�;"5�v�hyy9���Q@�*T���#� q�����V�O�f�����훆�n�@��������"��<I��e�ԔaхꙁS%�����q��gC���!��BހR��R���].Z��'����NS�˽��S����X���51��@��U�de=�����EFFb�2�)���������.�AڸriK�
J\�.�А��K�{�L=l&�%� �tn=zLU �s�YT�k�怐��*�/ �[V�I�P�#�?-��S�2�Q�f8			�^_ҫ��鱣q�M�8�m��aˍT�G�Fs  Bи8;;�&B�22�i��Tz��������� X�hwvpp�.��>ӷjhn���-�#�DṶb{w�<,�f���ph�ݍ�N��1W0�-�f.�ӹ�����v/���x��I~���g<�~n�9�#�CW����4��UK������UqkxE�U�u��ԭLM��\m� �
��+�iX��d��`�>H��K�`��?D4Uƈ��1���`���|�-f6�����e���!�'!�Nm�Em�|���~���3��@𼽗���칾�M�DN��U��2g(\r�L
x[f;	@���?��= 7*�s)i�::��knHYZQY�/�jL�L�M�7 xTTT�nv�=F���P��3c\��F].�ı�<"1}�͐�C�%q�U�sK�P�A]�?k��ܝ�X����?��#;���bm�w6&뫸��{�h��

/>~O46q��P�ݕ�f���-��T�;����3�D��T�*�rN�};��&�V��$˾˄��Y�p����DW�z�[WRRZ�=��t;��L|KK�������Y1����|>�ń�U���i`�Z?�Bu#t!�v�L���WI(���-/<��O55s�5���� ��XG@���p�ډ]���h2?\���˭
91޻�\ ��k߃Z��B�P>�98�HQ֋ET�>�r�W��y8N?	�(�ĖI�g�����W�gK���cBS�Z�z���,���l�^k��9B��u܌�7�>�={�=�u1/r���3k�Ua"��(�|��� ��''��yϚU�I>Ae�J�@y#<^?Vs����;B�=��&�NpX�I����nXoffv�kL��%0�(���6a[v>�a 9���yCf��E"�)��`7�f]�$�]�٦ŭ�֠Ya_��o�%'51��؊J� � #����nY&&&ݯ./�s�n=�h�t���<:<��a�r�_�v%�s###�<|C�^4d�u��6�Zzz�V��{ѴCx=TX-B�n�-�l5�T��u0a&XQ���yLNf�:�U��VA�WEd�HNps
7��Sm�P�[ʢU��gH
^�&�T[n��BLCm�n{�sZ���X�����RJ�@�Q^#�����B�쭢dD���_����x~��޾��N�U�f�'�X"k��B��Ԓ�?zNZ=��=��'&�� "��+ٍ�yѲǵ
Y��"^�0��������Swq&$Yd� ��)@���'�'!]H�����i�B!w�ݣT �僄Y�Np�������q�΀�X�J>B'��n��<4hO��˻M����Y3�Ft�gY��6f�HJ�����aZL�?b�7������C�&�: |�K����/���.��v�=��bD����
J���ǨIoz9�+�<سn=�Ye��r���lvlvZ�t�e�5�Z�O�����L�V�����]5�<а���p�&����	��R�X�޽{�sc]�Gkk��z����=]]����(���/P��D����?�d����db��J1� Xb8ɠ[Yщ����i�U��GZ|;�����?a�'��E�/�j�*��)s�������έ^>8d��X�m�����V����5�[wb��kk��YYY!�Dy���pe?�QQW9Mc;?�H��A�`����`������a�TS����C�P�ц���b��P9�,L ���S�=;�)�DwRy��ʻ'v��0wl���#PӽU1@)��"ؑ�7�#���K�s��K�.zz��d�>\L����ˍ
�V����tP��_u=�m�77�	����/��;g,[d|����и=(�w�����i�DN��)l8,���NM�;�<K,�nG84�V�Mn����-Je���A5�)�Q�׿��LNN�/|���no�g�2z9��}� DcYj}7:t�F ˿��q:;��� �<�n4�~=��|0� ���6�n�V��봰6��k�9k���4���\2Z�=|��Y:F>/�r�2J����T� o��%k	� G��MXweT���lƘ�@�V�C����C'o�!�u+�Kp@!�O�Q���2����m���]>�OXX�u�$������=8Ce���Р>+Q#F}��[l�C3�c�wo%~b+��O����L�"�v�<����:��/uA{�E����$���y_x��ꨗ����?Z���7;�bqk{�奥W����+�AN��U����j���[>\>��ȓf�K�}���Iw�����!=㶮�'-��s~��H�2�qv�Q&;f�9���A�*:��_��?�1��ۻ�+�>���3��A[�JbMi����8����Zb�Ű [�vOV>�jA26p���o�q� 9�Kk��핳�_�ĳ�g��uSܗ&�R7J�5�2�_���A���*�E�.?d��9�m��5�1rAΨ*�����ቭc�������;'v�ϓT����B3��"�S#��i�P����@n�����q
oNC��a�zdݕuk��ⴸ����z�V-�����}Z����!��.M��W���P8��dV⭩Ke��YCé��������ު	T���{�` ��`�d�k(V�|�"�2�c��o$��=E��o�=�X����U֮#����7�U�Z�}�Ү��$�~�M�T�f�������0����dts){�f�)a-���� W��"�����\W�����4�u�zu�;MMA�}��2������v��t��\�>#L�N�1�!Ԙp3��.���c_�*���P�aMbU���WTU%a�>��H���'�r��E�8���:bb�2�߱�1XM\��)@k�q�X����/��q��JC�8`��'R�󟣫]���I��>~��d�Л!�{�k��[;�����ˠt��(��H��x�K���	�\�<~�Gx4�A �\]>�ߥx`� �wT��@��Re�%���6.9��O��vx�����O��ʋ"�i��}��l�V�]/��$����]?���A >��޾��o`0��<���+���͍��w�$'�$�m�Be�_Y���/��,<�^��i�GY~FX���G��_;��-<З�k�~)�'���T��@Y-�2�Pk��)�Jt�	z��X��\�����wa��*��d�Y]�x�{������OK<m.] ��/#`u� x��ټ��7u�ఓ4��c����"o){�5X��a�v����yx��>�����4�b�_�{^Tt�����Jv�Ganx�CzF$��Q�6*3�X[�:Z1j���@��p���w>Ʈ@ȠE���f�z��s�	R�G�'�Ĳt�U�X�R�{&�ߛ��l����S�ј �_����!t;���y=t�p��j����x q ���ڵ���.��p�I�?;5���*�8&V,]��1X9|���q �c��p���R5C�#\Q;��L���Fn�qOv��i�<x��vAI`����G��� P�6�����N�i�A:�آ>1�v���h�Ž�e���^&''�9\8���~��QNǲ�{K��^w�ݼ���ތ\���>������m4�*F���4þ�I}ߢ��*%t��\����]�{��QJ!��G�5�d���o�'���n��)����>�z��R�����o}��K��5km�[^4��]Q�8w'���<r�����-�<���5�*�����*񓉿`{�x���}�v�������8�w�#C�`�g�����8�HUαM��s3)od�L�\z��ʓ����pF�T?��kn�v���"""�\�l���i��'Ŏ6����m77wZ4���j��=�\+����Tu�D:�Mks�.����giF�y�t�@�u���y%�S���M�	���_H�Mݙ��W�v��Pi*?M�ƞ�D�au�5Y'P��w��Br���X	������q�"�^/�u�~�9]N�BU����o�W�Pu@�C-�������5o˟XE��v=ټ�������^ǻ�qǢ�ϑukN����V���1ڢ��6�>�y��h����YKb�h��������R�+�Ŷ��j�#|�Rvm]��<f�0���}�*�����yA=��a#�2�7����������뿱���!җ��M����Cs^���z����T�]������,՜+l��C�y��D��!���300�@wܿ퇉���9,��L���m������'1BMH�l���]v�a�uB��Ύ�O�>f�����Ox���Ii���))zIu���pZ�, u�TH�Tz�j;�%%� ��^�Z�����?I�˝uLw���2՛��3	w�� ��w��y)�fo��Q�^�x�3��~�a���i��6['�#3�$��d�����̙^�<y-���4C�]��+��H�#J�N���)�9xpo&�]�=�N�Lo������
MMۧv���=��+����+r���K�$6��v��1V�a]ۈJ/L��j�6�G�;p5���C�c�c����&��%-iN�&GF~$�9��@`�s����orH))&��B��3�9�Ƴ���_*�~A�a�����8���m�N���X���7r��hIV�|�9�����u�U��m��M��ʡ�y�1U>�9�k�(P�/v��v��6���I�"Β��,U{�帏����0��K2h%��ma�{͎��M�x1 wz�d�6�*��Luh���)���yg�����L�*\���{� �efK���!��w�2E��X: 0��
-���'�����kHs�jD�WO��<)� �a�M�E��G7`��R�ߏ?�|�K?)dĹQ^OLU�&zU^��a�����=�a������/ճ���`��xq���b<?����TJn���Z	;��hp���C7R���G���8�M�zބ��w�~LM-�$P�������\���b��{@r(a�|����K��yŜ��#�U/C��Ƈ �$�O��	�lZ� )�ݖMt�v,e�03ҫK(�TOWO�GA�^��L���!ef��2���P0ˉ�@h=mnBL$�l��DC'f&�8��W�Oo�{s�W�����Z|g��3Z�A@�ec��]䕥2lоV�������8�Bm_ѐf�G�$�����Dc�����9WB������F�Xt[��ޓ8Ҋ�ɬ�{����L\�(a[mB#��;@�?~��=x�3�9�D��ȰJ�ղn��SA%�SM:]-�j��5��P���6X�n�U���Yv3W�,�3�k�sg���s�_�R��T�)���(�F�1�fB7�O֌YWT�r%���e�y���y���r�R�C���'���mG�>c8�[N��4�<�$����i�[�@e�Y?	�A�֮�q-��zM}.�RC+����k	Dcn��$Q#�����f��Բ��dMؿ9�(�v�K�̾*O3'5ѝ�K�'���NW���f��У.�YrYB����ܻ��{`.�+j�{�u��Mt�XX�r���t鑤͓�|��G��1���4�&�ߋ4JNpncd��j�p��@E��m��S�mo����ڦ���9{y�T���� � �'P�HF�f��=�a�'s�0cA�3��x��f���CRBܴAZ�AJ�Y󃰐Uԋ�)��÷��05�$�Ct�&x?&7�/��J�4F��rUc`2����ڭ�X���|���I��2�������,��vZ����׭3[�4⻂JL�&���h)��\?~��aۤ��iُ!�IX����L#R��H�F'�'���g����E���o~B��Zq�3��m~����C�����> ��������Ig�Hs̅7�Yt}Pa�-����1|���Le��������d�efp��C�����h��_��$Y��������V&Q�:��k�@�FN.i���C�$�޽���u��b�7�w��+��y���{��_�]D�Dcb¹-��^�M����0�h��y�$#2K_��13c��gX{A�Z����[հH,+�����7&����IL/��������H�W��J��1#Q>y������z�bE�����juW���4R2z
0z���R��ϿrH|Q��Ƣc���V�D7�XQ�]>�@����-�Z�a~s��1�[��7V[K
�#ď\5�����
!�{�L>T<h[Ĵn4��	����<|��Z���-��P�m>��C�'v�p�NJby(B�����!�B��L��b����p�`0�L"NQ�������t�^O���)��*�c��h.�V|�e������D[X��s6`O�.T � lۣ
U�ŭny�Oo�i�7D��v�:�옷(�������v��s�s,���c�6��ل ���x͝���$���[]���i&�Yn80�QD�Ɍ��	�~"�j2���HꙕC�����(�$�7?�X
@�1�b�[tr�n]	bq����l�t��BU��/�(Þ�c')¼�]����	�p�/t/_�L_�sn��T;L�^G�>Ļ��8R&&�gQ􅥺���6ޔC��ڞ�hd!��G6�F���(�h`��]4��@4_�YJ��ѿ��E��!��k���%~ q�Aa.F=�2R��6s����G�����ڷ՝S��L�!��Q
��'���9��r`�my�&��v��z��e�{��&R�.����
�7����&�޹Ô��=z���
46����@O�
��.Ԩ��l����"D�0�U<��w߷Y�����$�m	�a\q��QM����L��)x�O�`	��B!���ؓɤ�i�<�1�a�c˒��߅����t��;e/P	��.�c=�*H)�"��
jf���:�f�A�d)$&��L�m
��G�z�/{��۠�fy���=�6O���p��qH1:%�6|wV�77uQnL����"3Ӯ��NuAN�{W�x5�k��0�v�|O��꜊�PV
�su·�`�s�\�3�~�k��95�M�9�H��?,���wwY��%�'�@m_��b1=4���!����h��Xo��8#�~��� ^�
��`�jeG�0��h�/�) �FTD
d48�Y����dZn@|�m�_����A4�΄[�����5oNj�u=b��� 6�e� 蕰<W��73�3cU�	�0m�&Q#�(Pl��[s�����0c�J�n����v}<S�%vY�+�����󇣘3\�G���D8s�����D{��_+6-��=#zg  ��PN(�lԧjL}nX!�$�[^4Pw�d��²���3�ݾȡ�by����@Q�'[^@��A�,gXx������-Df��kk�P�/ac��k����Q�-�YW�l��->S�O
Rp�$�s���R��֏�"�*�A_�h��͌�&]G��57�8B�ω��v�z?�����@E��2z�P����Q����YZ�8$��n��ͫ��^BwYh��U9�y~0��K���	�,5?l��|�?�M���:�rTE$�6��Sv؊G��<g6llC+�K���W����de�Un,����@%~U��0���������/�Q�m�������:�O�?�b�b�O��rL�ｔX;f�|l�������@3��C�a����G堟��zhl/pfd6�LL@��V�\�d-Y����_fl�ņ��Q�yltX�Rֱv��le�$@>7���n��E�L]�Kגd���>8���^���؆^MN�(X����kW����B��5�B)Z�u[����4ڴ̴IHBj��2�$�1ej����&-ӪFj�֩���=gr�Ͻ�{�9�����]�������sLJ��"��4�|F�����gjh'�x5E��K0/��8A�`���,��!]��;�|q�+�7��<L�-�>�A�b�h��IZ:-ۭG+���u��0�D)��C�Q�&��+Zא�W}�okk����w�IAHi��B=�Y�X�����A�xMwq%I�2���o�$�*�$��A=ݪ	j�:#�l]T�'WQ�m����.x|<���L��������W�Cci�w��Kx�QbE��;�o��pJ1b+^I��{T�^���,���	��:�<A�yF��"��P��<$�eB�"X���=ɡ��ml<���'P�����Lh��il$Y�Tf�P
��C������{��Q�-q|��6�^��xR�c�]�&�W�lW��ũ![�����%8M���aE2N�Qf����ݺr$��OY׍��,V�(�h3��Ҕ��_@kTu��T�"��PW��T/j ��o�ow��֏z�T+�bZRK�C��#�gtY)���m������{����q�jެ&D��1
7i�Rى����9=�.�K�ܑg}�|��rf";l"��pz�P_��
=�����TÎ��WG)�K<���gp����ռ��H-k��ϺȚ�n�`FN�SY��ůۈj��8���>$��p�����׺��39H������5ԯ�/ V HRX2�t@���S�j�o:�~����P�-�҄�~��F�_5-~Gz�uF� �h5�2����눴/���Bj�6$�"��ދ�VP� *��-�r<����y�~P��<˝�d_��	)ӡ%^��[�7��Dˢ����͌DÄ�U6H��w<Rp �YD�h��
I Z���u=��I�
KZ�I�ۀ�Hĵ�wȀY�Q����h��R
���Kcd�HIIi�� `R�^Q��啄L���n�0�%5g��d���R>3z�`��8�Z&��+����"HD����gQ�n�n�!��e	�7�x��y�F��ӈ�s�:�܍q�ׅO�d�1>� ���<�!gK�͔C��#�u���0�!}�U�v��L�����>?Y��r��rVU��'d�4�ƌpc�­�C�]hY�o������#k���U�T�g����.q#��X��g~�s���2I�vm�!/��f�v�V�[H7D��n�k|~C��4~�jw~���ˆ�󝕽�2h	�ɀE	���GѢ���}�s��0�/u�F��L,\�J1X^7����Ul���C\��m�QUi�����tVR�͓�q�b����Lh�2��yl+R���ejBG�)0\Z�����Hҡ:Dg�״tݤ(�вaTVK�JН����A�O����<��0����0�����ܢA� o�L�,�����u���s+G͔;ۢ
��?�Pʋ������#Oٚ�$;C.���6L�zt{i�����y��˵(*|Ӕ��B�w ��+M���
�$UeG_���t�ؚ<�U�	쑠��*��� J=|Od��[�I��N_
_v\}Uf�`Lﮗ�2�ed��\X,Vo���փHi�ؕQxB\1 TA�#���;ri~��RZ�wv�c��NP��{��+���:�N�M��fn�Q1��0��MhMK
��O�Jn((�8k_�up��~��^���������f\�J��G@�re�L.	��17�2����hB���lP{�?8V ��bK��3��짼�Qt�(�V����dUݏ"�<2%P�'��%�73-n�C�W'�$�����0W��;�մ�tAXY`�R�>�
Xw��\�D>�+�:)ʊP��<�2+ `���ڐ]�#�����(9�
����q3��/�@EI��z��)eeh�	�a�ܢ	�Vâ�B��ىG6�K��(n*�0/�/*̣,"k��C�ޗ�����u[���ӔTӤ��>7�6�}i0%E�zSH�3� �f��Rs�]�_mG6���>N��**D92�4#rme��}lH�GV}���Ɂ� ��Q�V��s�$��~em0tHE�Yyx�9YLg�0k��z-������`��u�V�\l����p��s?���Ɣm��v<)�~}�Ŵ��st�@mKΝ����"�\�ʎ>S�4p�2م�����|�bA VuA�7��~��.��B_�B�w�T�����_2?�h�NY�ƪ)���[���_c��;?� n]�2pnm����V��LQA���3&3��f�͚��͹o����o���Y���ە�X��n�XQ�XP*�·xAx���e謮N �'�G��s����O�T.�Q�2V����++��ؑEu�	f���C� Ȕ��	��'d@n^2�* �U%fI&��M�Y��y鏏f���x�ѣm)=@ ��Y\�M�����g���?CA9R� �*Q�sA(��I��{�N��77����q����I���ć�D?H����$��)�h�D����Q%~!���C�Q�J������H�+�{h�� ��t�5ٔϫ�`Ƀ-S��ONN����*��B]<xkGD�jef}_��P��t��Qz�m(
D2v�>H��Ǹ�8�	6�7���3�$��(5m[����O��Z�����(����,�ݰ)*�����g^���е����>>�N1;@[/&�[C9\m�j���e�����S)f8Ah���)�w ��(�
Pz�}�ywC�k�Wu�	�������8!�0�������6��,e�b��\��.�|����g%���q*��B�R	��d�>��@VYoR�%V^��3�*��A�694�qA�MҼ�%���Z͍.�vq!�ڟl�P��e��J;	��\pLo
6��6���u�P�����I��@�w�Ϯ��/˛�=�SD����Pq�z��G��{����ܷ-h���s!5"�����9�a��?�rz�c�@8ňn�����7j�ɵ�ؔ �[��E��.t�wf���Ҹt��j�����f�I���1�0�{ ��:Kɨ�bS'�p2��o*uV�D����&j�����t�{��v���m�Ƈ09.Al�ٽ����&��":n���\�n����J}N���GMF^��@��!ڟ�w" bG�;�H���|E�{��k�D0?Rc�����^C�͡K�%��:��yg''&��)7c�4��#�J���R�Y�~���g���oŖ|��� b(د����Ǭ����*r����p͚���;O�2��,y �R���(���?�b�9J�2�e�#�!Hk�2��~��^�V:�����{�;�>?K+Π������Ȁa����	�*JO����_����h=���g9�mU�����a�7O�Y��+E	"I]"����ڡ���
n�k2�����V$K����6`o�״7�^�X��k�"��Ҏ��S�9nn�q*u��ɱUXl�)��Ԅ }����u��>���vc�
[�繞?+	i���iu<�^�t�ڄ��l=�գ͏��G)�r�ҿ�tz_U�l��~�Gř
:��5̧p�$���� �\��НR�}��@��j�l�Nj=�V�iR�i�3?j���B��Ղ�6~��F�ی� �m��q���0�3h=�qĎ>���w���L���Ec��ؙNl�i��ψ5IL�ep��	h�U�|�0+Xw��
;�1�C���$�����Ԫ�`�A^d=*���5�e��~�T���b˒�~�)g�7M��ݔ�p{g��X%�R}�DMg��c�j��^t�x���m��J�.�Z��=��/��J$N�<�k��"e��V��^8ß��&��e�V]-��EcX9u{}��7ى�ѷd���aJbD�ʏ���_A�����	Ʊ!K=��u�or�n20�7�Z�(	�����1@JR�&0�������\A�����P�vT�X�B?�<u�q��}�U7�x|D��g�����)t;dr!5d�&�<U���^z��)�"n�Y��)�5�9��l�+����k��P=$�����)!/�U�`���-��'Wnk)��|��p��+L�8��:\�0hw)�$�φ��9�=�� ��T_�����Q�<�%��r���T�����9D����p�\�{֕iL�t�V�&��rT4��[li܂�<гڷߖ<j�N�+�����q����N�4�ݞZF#���$ vTe�B��~Vx�d�$t��H�-�Ub�
�Q����M��t!�����'̘���f%�4�s:���M���7Ц���^��4G��؎X���Jk��$�ۃ���m�:�s[��쓂�ؤUp4��No{y|�R��,O�P�\��`�S*�&[�%㏻f'�咜��^4�=A���A,9*��*f	���M[˹ҡ���3�.0J�H*�ҙJ{O��.�6��6�^�d�������k3�img��˺����y��?�,vBx
����BV�˽E�A}ׇ��+�O�#=t
~$��tIt���l�+����ꦻhX�_;�����Sߐ߂Z�1Ur��x0@߾$���8��υdU�%��a�D��F�K0���vvT���ԝ�g4HDr��s�y6��G��uUUT9�y��KD�\�S&wmg�� �E�4'�bJ��}��'#�P������<�5����3"?�9�x�Y����xv'�N*���Я�?F��m���T妌��\�:� ؅�)N�%��� ����xň��\�āj�q��u�B�Y �jT���:�9ъ�e�~��V�T��Ր�"�p���ŖVn���I�F���I������9℺m�U���k+i=�� Ќ_��諬Q���Y]�����9��L�,`>�d�y_�e���|T�Hd �x�z4g��@F~b ��"��OvĖ����Q��s���L �e���8��F?q���{'4Y3�r �?�#~�/�`�N~��(��Ӌ`@Π_�)��#ܬ�
Y�o������R�E
��Ub]p��$�Ѧ@iB��\��P�sb e���m�0!��5{!�-S?��81���pU|~��H��UW�-S/�?�4��u���\]����k������5�x⯸pz7�������>����O]g��Z���V�{����GP	��z(��u�Q#��ٔ��4�/�S;-p�3٥'w���u��	P�:�{.U���f�&��=��	ƈF���]�%]�l1~3�'�]����6�c�����>�޳��@ˍ�q�x��b�;��E�Ae�25ի�=
�ՙυ�A�0�p�%z�`�����5ď1�P���z�'�ۈ����i=�.��㫫��nU}*���e����BMP�������4��:��c@��=Y��A6&��e�H1\��p�w;����٥!+�#GЅ�]O(�8w��@($�8��,��@��xָ�X���2)3�:q*I&������h3�W���Gpr#��4n�=����A럂�+��ۜ�9���lquI���,n���M!w��8�>�;��/��sSx	�uKD�h�WV���hT��E!�\$ӥ|�^ऺ��RՃ|����,�d���ɾ^<��{����4'5��)����J)=Z�P�]8�O�����{�İ�x�w���m%�<���Ҭu��Q���TYF'��;�*>0rs�fM,M�������i�����>�ǹ+	�������@=�lh30h�A믛��\ŖӋw��r�����D6ȡHL6`�e��p�1��Lߥ$ӽp����3���@����U��>��1�8����g =�>Z�u�D^]HVJ�"GsL����C�	IF�e��e����XP t�k�4?J���K�8)]˰���#�T6����ޯ�wm۸W��NQ�v�,���?���ܳ�9����)%�n�OA��{�8���eI�'�ڧ�I`e�@S��O>�e�)͎�%i��@���^�>�p�
����9��~ھ��:�z^X4��3�#u��o�C>����� !U.����7�^oRݢ�M払kH~t���+�d5��! 5:<1����z�!�U�U�:l�yM�������`[�!l}�^�DE��,YZ���J�󃛹����0'���ك�O~sx-J��C&@d�a�O�G��`�p&�R}��Q���Z[��7����ꝫ��[��ִ�w��y����w�]��Eb��B��#� v!�,S�����¤r� 9��%{e`�hˋ����K��:�)BfK��-�M���t��9+94?�17eبu��-�uq�gn9��7��ng噴�}��v
;��[��=r��Rrު>ǌ%��E4V���n��u�t�=F�A��R/�ܝ
s��
,	�i���#f�9[��ھ_��z�e��5Gu����6�#m��L=�����H�
Ğ��F�����[g�Jg�i7�T��p�p�VkK�&��j��ߴ���#ძXgO<q��*a�&	�52���jæ�����˔����4x�H������p��K�z��=Б�<�<�7�������>#�X��%W��5L\��:��UK������ȗ+2��r�`�"��"���U�~��p�ls?�5�Ͻ�{�����ɓ� ����q�3p�}z��H��Ƣ%�k�ƇW���_0F�؋��LCټn��<�K��\�����
ŁwEFH�F�2�J�P�c���xv�7f�X,�f���eMKbT����;�����+F��D��#Y�%��t�m=����7k�ȥS���y�)5̧�>�Th��}�ޟ���P����O�7����� �m�ОJj���q�y�ql�ǭXҺ��K�N�����V�Uu���*F o�#j!��4>�{'Wb�V/|U���I�y5�+_ݨ�E_� �B�b�}w�ˤg_��>�藏)�����ΫV��J�>��\����V�	|��Y(��ִ��񴞕=H�����r��ִ����6�&Y:#o�X��5�z���s�n&PM|�E��p�R�yb?g�2A��4$��1\$�AW��\�:���{7G�wU�(V��=*�D���\����@T��IX-����	B��2^q	Cf�A8R�8��"qj�����|�2�!AAi�	�S�N�E����O��0�s�k��!L���4��B����LOW9�]��<�j��)�^핍<5Z`B_��H(=�2�î:˧ǎ���JF�m���u�қ=	��};���Px��d�]��X�q "H1��%'+C�5�{2o���fHY:
��S���u��X�����a�Z�)�/	,t����݂?����/q�J�T��X^��듑7CQ:t���#��y�S�
�M6�b�l|1�w�9Ã�ާ��tI�A�U�ꈂ�F�3e�3z_N �W�`V�·��'��3n�{�}v�&���C44 ��#��P�vW�
d���˽x�����5�z��Ͻ��,@���7�X:����J�*u"p�S�t��!�Mk����Xx����%S����X���d���`I̓��ȉŖ��t?����o�J�:<��2.`=�V�����|�ҊsHd�p�� �kv��=��q�冊r�Q
�V���Q�/y
�o�O�	��k���Z��H����C]>u�s'�0�J,���l���,v�
�u�J���Q�=^ڴ(�O]�M��:����+�0y~��2����Y�$��6G���aH4Me����z�V{����3�u?���܌8q�����J�"������⦐�G�׾�G��5�..���eǷ��6�w_ǒn�v;�����u[��`��'d�m\-��sE,h�E�Y�rB��'��=_���@$R�l�mpnt��Ulil�؈���ν�H�/���	��̴o�=16�&������df�ңµ��ҋV�#坨�n�UK���x�����+RXn�j��a���q�Q�0-*�����.�f����h0�K*[�
��ŷ:&z>%w�7�-:G�J=Ƈi\��.~���"
A��8�vJc�]u�uc�RAn�c�V��K3��9��B���ߐ��{���ϴg��<��u��Tk�\چ��q���VǕ^e�5�/�Q�����K�e���2���^��s{��"M�p�,sO͚I}C/�2	%=�o�t3xn|D�u�/�ۯ�>X�|���g4m#b\sL'�\C�IeG_Z���NYm�Y;��������J����e�X����� D��w�e�g N���V�X���^��ye�;g���Pw~}��j�R���R�(��-n�H�"����J���π������G��CD���2@�|p�1��Y��׋i5'�tfH��r��֡:ē���x=w5�	2���^a��q����
\o�
ը(�4����ȅ����
��u*�"�o��!�\��򛁫r�࿅?�T�uF�W&�ͪ�7IL����n����`/d��9p��L�KS����$F(�U���@�6�`�1�iJ�Th0+�z�n��3@~����K�=�ߊOԬ'/g�& ��B"f��|Hݿ�7aZO[.f"���h[y��lB�x	)�ꔠË���E:�X };�X�����s�Tlu\�>����b���<2��L�[��9��$�,s��=!�� �HR);q����ؑMe时ܭl��0qy���j��������wHVAC�;�*��3��UF_�3�����>�����s��$�j6�T�죑�"�$�A��Q������2>.R�٤�{пI�[#��B�Y����V0/�v���nCۉ�AB����� /%;�}[*�BkA`�e�+�NPS_�j�RcA���r���WNK@<�'I�!Зo�N_SSͺ�tu���&���@�Ȍ�vdnJc��^����_��?�[d�,�y]>�ħO6M�2Ȉ��Wʛ�F�X�_f.�@$�o��x�}<��0���󲀤.uI�"��/�p{|n��2�%$�����S*'��$G�'��s����%��aNfk�-�4�=.P�'�j�F��!7��{ŪĞ`�2�7e����~r�a��!5g��=U�Lm$"<}<�=2̼�=��d�$Њ-���9b;�{D'���γL��I4MҊO�ۜi�V�A��&ܱ�C���-��U�5�%�
�vH��W��
$�����F@���7}0#����`� `޵*�C"*F�:���.[$We���w�#œо/uu��<��B����t���	������=�~��@��%9F\��<Ͽ�����Iap��E��8M��,s�w9u���_ܠ��$�A˰Z׀ŐI�L݅e�9���ݳ���N4E�+<�{,��k�jͤ���'iޖ��!��'*D��y	a"���H̯q�0X��"�|�+��q��Yǌ���	���G�<�$d����mk�����?�Ѹ���a5{8�\�)if���k�_Nѵh�:PF6��w^�<�(��Gk!���Ʋ�8��܆������b~�x䢚L�D���Q�r�P|j��:q��kBu ��з��s���b�Ě۟��&���)�MB�Uvㄝ���/�S�a�����@`�j`e�T�M9� C�Jp̼�Y��PS$\�A&�j|b����Z[��+Ig�O��`���B��s���|.N�
�h��z����S�h��Ye�i1��?�/�N��Q�^j�b��딖�ִ���GY�^���3�*��1a�Fp��: �C�bA����-0��Q9iuZΝܐ��2ޑ���<�=���q�jS����V"��	����=���F1�^�+��W'��ݥx��|����Q��@7X�W�v���Z&DV\�J��kr��5ή�e�4�n������n���]j2�����}�I츔����G�3��	<�=ئ>�(�zT7/�jfs��u��ߦu(������<u���bľ
C����h� ]iR|>��Z�b E��%9�M�,l	}VH�>?pRk��`}7�g���`��T�ˏ#���2c�j�r�
[���{�Z��b��>rFM��4��)�V�t���,��Q'��}�� �'X8����2d����}87C$��1��h�L���f"=�Ey)\L��QlyL����s̓��f�]��Y��c��o}���
��l����r��l�-�|���agN�%�J���Y��֒�w�WL"�ʄ���C�-#R1\s�����������ak�Z����xĊ]�X��pe��2O���B;�\L��	��7��v]ǶR�A�Nh�qB�S�g9���D�*�w$<PO�+q}������x��S�c�N^7Y!L?�Ɗ�kn�q}��se��N_l�>��$�P[=�]?$��b���##z07�,�#��d�]�ڜ�W��j2�}�k���;ac󐧴\ ���5��R�����PË�*�OM��#��i'��:��}����X�ܛj@����W�)��%ղ
?U?	_�*/D��}��ed�&n��Y��4mEۚ�˗WbI�I&N�ԇ�$Ӕ�L���B:7���ZBab>��������%�4�*e/������q'��[V��?G��,�y���}�*)���v�l���MC�t�ܶ{M"m��H˰�mc'����O�ұG4���ٖ���f��A��@�+A�p��#���C�$K&�}j[��|�4	g�O���z�,O�s��N�Qz�=u/\�b����=�w��P��4��g�g7���Qz�j�8n�	ͻ�3��$zȅ̺U|f�j�X�~X���'3���e�}>"��u�#4�Y�f��㋴�/_��r3�e�w?��aa���1SY,w|-V�[R^S-�lPP������j݊GVI���S�R��j�͉e13v�r�:;��4�71�,�`fCO1��C[��2I���������mBoa�m���R��Bu��f1/��C�+!P�����aA)����!������k���G.�
_���~����0���!�k�|܀+n�|�,��r*���]u���W����z?����C�0��ۙ)l�X�c��P[KK+�ZlB�9i��yIG�������'v�2�n�2����D��y�9c��Ea��S�3�[d���5��Tמ�ձmd]�OϬr���̨^���V]'�Z�t���%&�EEE�w��=-%e��u��L.^\2�����n��W�o?7�}�Q�����L!v��7 n���S]��Ȕm�I��}��~�}�F��b����5��JO�J���i�Yd�`<мY�36���]aWߡ,?̀R��}{��y��7;r�K#m���}ylfX3;�(nɯ�� ��ҹ
[��I��~�c�������MSRR�;ܽ[����N����7�_3��]�IE�j���
r��@׫)���qx��B,Ľw��w�RO)F�ыJ�1��͛�ҡ,1WA��t����C������T����~�	��p��2g���-4��ؕ7Q��~W�=��|�Z뗳 \l���,E�sد��<��f�R�:;!Z̧�'VJ��Ě$Vfmո
�j&��`��5��1|�T����d�S��,��~��|o����m�qh�����Q�θsh����ǅ��/wk7�w�*��`"K��SE����3*Ȫv �ʧ��Ыx��p��㨻b��5�Fj*�=��-(��e>��ic�(��SfQ���0�m�q��7�&�L���M��\~w�V͓����~>�g���`2^����냅s��7�rX�1�P�h�9����+?��^  ��7��L�N�5^�e}�@��P[�}7ke�G�{/���~p���^#�W{��U�����-��a����(�iZLy�7�a�o�Pg�i�xr���5,���=�ͭ��J��v�(�ybL����E�?-�I���Օe�a�b?	�l��у��3��`FUK��9Tّ-��Fe�[~f-�5gtCVT��,���h����)�3iQ������L��=9EZ���	h��XO�1(/<j�n��/n�r�-�r��8f2��bL�'���}�'K�vm��E�ڵ��Ìyc��t1��;i,�~�� E��d:�2�����`+�H�m�X�7�n��a�T���p�yr�z?��Xr-p�]��$w�aB���U�9�a�ǖ�� �duw��x���<<CU0��e�3��O?�Q���$`�⅚r	RoI�F�#�D�v9YVd*D}��❕��T�Q�������_�7�6��^�8u�`ۻ.N�I���l�aΫ�}��3]�|b�3�F<BuVm_�����(R�ܳ�	`KA��U��@�XL4M0v�h�/����jUԏ�&e���6�������/�~���"VR7��H��dt����uƪU*���rm8�9P��}�m̛x�Y	r�9�O�R�,��7b�7����:���ۗ��|���dm�F��>���{�P.㸥�+�`v�3z6)*�>v�ݭ�=K,3����:���傉NY��s|TK�G���y+JR~�%M�6ZC�뗴�1z�5�0s�7�r%��7��>b��Ev�b	𷫩3�D��7�mhZ��$��&E�%�B� ��,Fx���ђ3�M$�p,�PN3]�h�b(c��V��L����։�s1�Χȵ���}�^�*JNE9KϝF��.lM�|�2g��`���;p�@y�B����@��G,w΂!���V�ny��(������CC��T��	#O�8&UN��:s��Z��'�;l�R�1�Yv3�2,i����Ab����PB}La��$����̆��Ia
��v�Al�߼6��)�u�3�%�_";�\�$��\F��G�V���,��>rєo�$�iҽ����j#܃�� S�1�/;Ny�d;f�e�f&�N0n�	�������/�V��ߧ��͈�����T������������].G﮷Q���0��f�w��i�v�r�B:��oC̶��i9}nS��;o#�0k�$Y�L��%H"�׈D�Ȣ������#��b�=���<���h���'I����3�d��ޠ$�&r0�L��M��u�g�����9?~��Jp��(7b!e��N���EK����T����)�V���Z�&�](^��S߳����>���@9�f�:�D,[�a<�Ŭ�B/�ٶ�L�J��s�=���ց�R��5�3�7�Dh�-ǲ}��է_���O�Z>Q�AQ����lzī���s���̨*���u�'���5gF��7��$��Vl0bs`����Z�bK�JtԜb�(�x1�[7t���<`ȟ�!��c�KMƼ�����sg�%�9o����C���iy}|ӫ�Ҩ��Bk��lIq1�jr��N�I���%�������ғ�eu	�ԐKΝ�靤���g�H��7�9#�̮2	F�S�hX,`�CȞ,�g��U
g��=EqhX���c���r����|�Kq��Xjuuu�� �(x�� �54ߪ���{Y8�{���d���j���;9�D_p{U�
�o�4d�x���ؼW��g��@�`�dC�P�PcqK�ρ�w�ಊ�����t�v�/���R��xl�$�xmQy�'���C�r
=�=�*�	Y�Q����f�� Π�w�N[�Pc�^��$�S��MWՆշ����7��o�::
7�r0�6	���ˊV!��(/ 5n�<����R��.���D�ކ��jY݃�������\P�I&!Zq/F�}�����҈s�,����g��e�~g{��v�ўu����sy�qm06\�Nl��.�@�~�^F5ߏ����I��H`%d�{��qnh8�`��=J�v�Q���o��gx'MQ^�k#�������g���S"/Ci�K�i�|Ts���D���f��%r�Ѕq��򝮦�,LhW��֨G/-�ֲ5����J؁#�!^��o ALy�W���l�����ó��Hf5�?�BU� ���60�[�����i%�N�l4�%����U���xh"��ǎ�|\����I�T��.��1�?H+Σ�cVvUG߹�9�@����=��z��0�����<9ZKDn�9�S7��>�ju>�Z;?pӦMe��Y�<��0��P�0�(������Ͱ��W<�Jvϩ
���oFo,��jD���`����r���2F�[gVHPP�KCU����z?�m�f�=5M�z{�z`AĻN�u����v��{d�n���&Ű���+lAv�S:��y%��(檻�D��@���B��BC�`'x���:� @����v� �^UX8�+�-�#��ذA]f�O�}��O��+��NO[HB,Snx�y]����v��E����c��z��!o\̼�Wv/�=�Bne<���HDzNq�����N�\�E������.�����S����7�[�])[)b���s܏�j~�Q/��Y9��3��9�~������XnKNr��>I�����<K����l���t�b���$-�I����
_���YJ�RǅF	���AdD����Q����m��W Y+� !:������~Ո���Ndɱ�]j�̬ғ��M��{l���-�?���L���jT���iV�QyW�����o��9�~�魉��!j�҈pOU�{c0)�-���<�ɓ'����Z9z���́���r,��\��ķ�zF�-az�Gd#����}�.�rd�9�S�N���W�;����/��x0z�YH�SBv~����	���@��*^� P��\���u�>�����#�:���j��vg��1����J�.�T*0>n�EI�����	�ռ���?�2�J\;w��6nc�{V�������p��1�v��1+f��$�"��&(�t��g��u�)d�1�i��`��SI��0?�Jl0��>/��Ea� ���x�?�m�(��L�|�K�)���{V=�t\�U��W'a;�P:Hݹ�O��������&F㮢Y�;�;�� 8D�e{����Z��j*��Uzpo��*%�}޴I` Ǘ�����=)t�y�BU��O��9�p���B�~��/�=�=�Oڟ�������[O�L��l0����q�wj���1�~	���:����lx��������;�����ŗ�s��d�O��_�1(JIB��b�O���c����M���V��n�l��Ґ�I!��4͊��Ag#�u�׻�)G]I3Mb�r��Ǽ���]��)��-�����龙�E�OY	t���?�k~����
��[����^��%�Ǭ�\jr%ֶ�؄m��'sB�П�{��18����'��*6��w���]��:D�	I�3rW�X��m��s����d����V�P����斺s^i��aC���ȹ��/w{T�t+�Q9)��¸��~�쿩��8�8q��uS$�yO^�9�D��)�׻n�C!�&��l�m��o}l*=��Q��p���)9��Dz'w5�x�ɘ�Fv��,�0M�zZmx��o���ۢ�x5A���o�Q����?�Y$Q҄��͓���\n�e�߲�w�e������DF� �C���WSL�y����~�o��o碰޷l�l����������]����A&��%�*���S�K���fQ��.���ŦMȕ�R�;��>�p����w+F3����k�B�"iD ׏�d��U�w���W�y���E�~ӝu+�X'�#;�R��/�OR,S��\�T[��Y �S�~�?!��I�RX>��a��D���D����@UR��+��a����k��粅}ļm_�yh<R2�Y�%�N���_�;�n�l�߸��Ŋ�w<+�u�b���W�>��ۏ�c�^��kyNY�9��ԿÚP�\mX��`��?���^&zԮ�'���]�Ʒi��_�&���r	���Z�� �ɈW��٪���߭���&_o�rd�z$<	���1+3�Nc�v�{��9)	�)���ǃ�g([hs��Z�k��x�ӏkm_���7���m��|��v{5�UP����:4��yy]"�pEx;�X�Py��rC���bNi�h��<&�<�D�?�.��;|%��_��{8r��/ZY[ �t�{��Y�7�jk�[NL��W��eDC�>E��YƟ(
�Y����z��?��ť�v}�ȿ���*X������3��hm%]��/�%`�P��$��|1&D��(������"j�V�)y�m/t���^��:�����7��g	j�֙e�4�Ջ2E�������{��H�1��\K׶�^1����+a�� �f �����|��5�~Śߑ������#1.����[�� x R���]���ъ
��w����_q�\��aٛD0��ړ�3f��@_�b�җ�  �:�W<����աg<fq�|F�7a�勲� I�pX���*6��T�?Dn�AȌ���
��g�/�}KPF�$p�o|�9�EX�U �l�L�&���o&��be̍v��
�r��!}�C�tެ��Y�n�i���w_�����2�c�htRu�D�\��o��/�"]�	_�Ԗ{��GA\��Ca��� ��m�'ߙ*������`3�)DWl�lR�0�}z��b�����e�1 �Mn�?m�gF\!��_`�or����5L�����_�7��zFq�ػ-�E�:rQ�|1R7Y�T2�}����a>�������������~�z<v/Ť��+Uk�C��2��?Д\d>���v��i�$�"}]�n���S7k)����%��c�ʡ�Aw�o`�*.aF�Тܒ�X|��O��޷�,(��-p#?AϚ�*������!�_�^?�x�#n a�5m��<x�Zk�	kň����I&�&&&w�v�I&�f��)�&��}ͅo>~�?wڤci��h&[�6���HL,�����9^�A�ŝ6��ًo�Ǜh��ęg�.�_�����	U��J�v|92���3�ׯ_��q���N�Yصk��携�젧9�ǝ��_��	J�`6ٟDb
b� 	MdK�YZ�ZH�~LAY�!7��A`�b
��wuw;6/;wF������\+�P*|��Mu��իW?zt�j))���� W=b�Zz��H�������BY�Q����~�z�W;��u�T^���3?>UY�n���#�j��9&���ĵ�x���,j=�}̼	�7p� <BF.ZF���+@D� nW��#G4�ϟ�!?D����(<&�`�j�vjń�!���^������ݴu��Cd���|����KUpo�%g.W��n8f,9�a�{��W���ٟ�?�7�Z����CF� Ba�q����a�j���c$�k���I&'�Y�}L��,��O��8X�����SU��T/���s0w��p8E���ÙX�f�+��ơ(i=��fFuͅ�r�vvz��l9''�qv��UQ�"��Cd��0�_Qq��>��S��w����,�NF�z�m-f�|��e؆5�KHNF���}M�w��������������+�8�gddd^N{�z�LA?���ǢSN`�:���+������zz��S�ڝ���ݻ�~ih��w����I^~�]���a�Vo��DÄ7����Y)x�y5�>��NQ�b���?���ԥ��RE�q��m韃��=E2E�gյ?U��!�R���Y9:"C�����n�޺.C~����J��'zzz�L�_o�:�W���u����P��[o.��AS�K�'�;fD�݋�o��o������M���%��7��r�M��v���rؾ�1W-��v���}x�tYyy�M**내V��*|���W��?��-<����s�����g()��� ��S�f�!��$%������,�]!`+�ֱ����#UW�仞?ZZ{��ZC�h|��]s*9��oCC3��h�3����#_��� ���%�� 1%d�)����ǖm'^C���O脻��̥�+�H��;qv��H@Ӥw�dH�Z�
q	��p����E�G:UUA}3)��͛W'�|ӑ�-k��uކ�̥8x����;��j*���Z5�����0��R\R����>�c��ݬ7���6o^�Ve�sx����������L��E�I�C���ȃb�a13���Qp{a�O�_�[�)/�Ri}{�7�Α����7
[7k��&�F���iО2O\s��h���1�{�\���4�$�s��*����rZ-�����T/z�4$�b/��8U§�ԛ�a������C_Kܟ\���k$��q�R1�B��̮�b�L{�C�a���ޕ)<�od�`|��r�o�:�Z�[[��Ɲ�\H���w�)Vj}sm�&e�[�+������&ih��xx�`vY��nF�陳6u��: $Puʱ��[�{�/Qs7�g�k����Kg�����U@	��i�f�����F������>�&�y��	��� ׻�^W��h���Y#���ط�0�?4t�`��g���̮�)��N���7�����>�L?���n�A�N}��b{��g#�:�����9ͯ��V�GD��n�c&+U^^������#��<��1�W]��^��/�� /L���K2��ӂ,~'�� �J�l�@~��W����1ⶋ�9�Mv <������$�e8I�罸ZM�'/��6��TeuKK���L߅�ՓQ���Z����n��pk�����>��{��f��<$�U�d��kS��W����.c����O��2�m�+a��ۯG������1�G�3=y�a��C��={�Ν��Ŕ���w�`<����W���\x��	3V�V7X��V���[��}�#���>SB]f�S�?����EA���p����	��M���a�AFL��D��U�-o����
�7x��1kB{[0�����U�of C9�w���?��;@7���ܞ+��������Ϸ� V՚Ɩ��ucI�<[	�0 HB�����EQ)$��>�Dqyp�-1Y�g��ћ���#��[mS� T��z�S�]sYB���H�M]�����c��án��qWuE�R�JYs)k�
)BTD�Dd_�eƌ\-�W*���(�2H%Q��B��fb,��9d�u����s�~��u�}>s��>���z���C�J��i�?[��QϬ��^J���,.a=�MӚ�lz� �ނ=nhI���~Q2eE�+8�~ګ~�B����R�˰��=�!VIB��Tq�M�d�D2�Ǭg8[����9yKp2?J �h�Q�����r2ژ��:��n�v���+5\����j+(����m�!єa�ߝn ڐ���Uw�ݾ�Z%�1t�'����랢[�����c��ڋ<{�>�QɐE�<6�jX��d+;;��?�
(3m�K�x����\~��M���PVM����W�5�doyvxk�����R�Ԉ3��[:�1.��%y�5.��oW�	E�Ay���7���W��}~�`~�;7k����!\��!	jQW�|�#G���D2��ܣ� R���Z@�h�|	������:�t���y�s��y�X��%WRJ�p��9�9��+H�K�ȺߐuϝS��"	�'� �����<|��p�Ǉ�R���Q�H.�߇��<u0X��C��&@I�
5=Hm��jH��Q[���/�AF���|e��>�V�9Y���:1�3'�Ո��0���¬�AR�++���-PJm��<���F>d،��B��_���Ă_��-#��t��*.�!�L ڞ�0����;���2i��%��m���-*��r	���?�i�RQ
�H\�pLlS�ϑn�q��ź��1rEL�H@��j��������ɽ�2;i?��8{��:nq�~v��=�����{��a��q`��&q�����4��O�������bf�vxJ�R��]OŶ��,��4B>r�:ɤ�KO�$���q��̞���z�� �IT��7o�J"���4ӫ��2Jg���0@?w�T����J�*��.%�L &fc+=� x����Hi+�4�o�L������N��sX@�1���<Z�����2��S����B�ɻY�F�8��s[>��W�[�~5�{j�w��$>���I�ܰo|�ج�rF��[��[�P�Dq��������*��e��/�XS��D/N��B]��t���+�D\{�9Y�W�t2�t��Ą��1}+W	�k����mఏ�V���.�n���N�h�XgonffY:���69��FMwoj�-ܳ��O��Jۯ
Mo u=�<P�p��Gy���i&�B+w�*���U6_8�1n��U���8@���O�[o d����䪵e�ּ^`Bn�=G�s��Ӽ�eQgY��6a���aV@���sxj@��w.�+�G���������9b_��dO���������ڵ�>}�5=<7K ׳�U�ZH����� �D+��FDx\��G�X���S���9-H�gʊW/��#�#˦&�-r.oo��W��.ʹ��5H�
�7�����S#����>?�S[�v��G�v�r����&��&���	+Fa��=R� r4v�J�jjY �'Y��q�&�UB]��л�H/'D6����9�-6i�~I���n��L��\z��Ț���鑊ѡfi����.�1��,��j	X�be�;nWEHj%���_7���K=-�=�ȡ%۶:l�]������[G��sf�J���BCP�F��^�Mi��+[���Ç������!�~��3&�<J����	lY!az����:�u��GJ(�᷐Sկ<V
z�A����>���EhKA
p&�E�L��`���j��

�v���(�:t
�ŝ����+�
1���:�D�م�V&!h�џ LO��v�X^Ҳ�p$ 3���Syw�7���n�)�LZK谂���b �+..�V�'Towǃ�p$��yQV�X�*p�VK�R�.��pZ4
��IW��2}�U�k���ԀOw7�G�rF�'Z^pBR��O�y�
�T�#�ϝ��Q-ZO;��|8'��S!���<҇h���{[�"aI�^LB�]r^$��e���.G$�g4��ҁU#���!��ȂY�õ<�h�J�QCԔ��	�X����u���y��=*��G\;���h��j~����gϟ 8�D���ocb���[�1�W�čMM��)�xR��]��6�U?�@P͇Bl.0с]_�%�~��&��Z=E�3O:��Ԯ��cG�X�2Oػu���lq��xOXN�cJ��� ���f��J>l���ڐU��9�:{n�]�\�d�I���������WdP��Փv�=(��X�Xh��ћ:ɂ��gf�^Ļ���]DVAU�9@� (��<�>{&���o�$$$�m�vT�p\t��o�:񇹳P�����N3�>lHXTT4[q�'��"���%��@��M�w�0�T��S;�B�U!6 `j�p<�"�V����JN����r
�u!������9b��O�e[C��������p��֬Y3
>@2tu�����e�����0>��˔.G�^����c����Om�<�o���A!S�b����/6�:HVx�:=]���slo��7y(r?�,6j96Y� 	�d��~�	���#��=���Q�۟�GsJ�i�h;��>�[K~��V	��iW�.\��B��mn[\7=�:���{-ÔV����85�yGuu���8�J�N�"2J�4;��CN���@�«�t��3��V\㜅�ߤ���'�u�>N!ԁ�=o9
\��h��z�Y#1C�YI�ɨ�t�5��r(��e1&4���쨌����	o�!�d����䗆�DP"�h4�B��o�Qh{�GT�=1Hu��] r(�I33�ލ�������|���ݗ����ñG��ө����f���S���;�0m���}����7;C�t~�-|ں�rnĖ210M�mr��Sy�k����ݮ�ɨ��Դy�}Y�[Z��ft����\�*}�_w���K���q�}��'�WT-�4��a<�Z�]�q��<���%�J\�}3�؟=��]̧�s
T9���'�
�s�;ʄRÆ���Nz6� w��$E�N<�;���(*�f�*V��yAGK�c�l��*j�uΒ�ι��5��u���%
(�]V:[�x>��hkk�8'\SXQ_�v�=N5�������.�z#�*�fN�%ⴷ����C�r��v���������eio��?^Gmz�}�92ύqK���^~u�ho��hgbj�?���izf��_�}���P���d��9=�CY9����M �j���mV�;.�(�`��|��g�5T�ˏ�l�{ǼQS�"J�����ㅆ�ZrR�#iw����Us�cG{��]*~|@�`��PJ���:���F�E9�C�&�uޅ(��VQ#tۗt�V9�Z�)�\��C���̷��4�͔	���gCC%�L��c����E����`Mg��@�ț//��O����"�7P��b#��N�ww�JKi<����@n��̞B�A�ٻ4��W.��n��"���a�͐_��9���C��C�W[�K"�|���R�� -U 3{�)����1#����ֶ�^��{n�B��:�9Iu��|�ѵ*������_�]48�-|��AXuﻍ�l��ɾ'\�+��#`���ùdr�����ul��_{Fu}�蠬�0:����X�����dv{3���d!��63��|��ݳ��t���_�	�@X
G�8�5����� b2��/��?� ���YYaD�zѮq�̾Ч#��m�S���+_��[h�+\)2�[y��Cһo[�=$��{	����?����T��܄9���]�b|<{�_C�����)W}tm�Q�w�����rZ\%ַo߬,,�T��x�;]���)�*{�Fɭ�UHJU���-|t���Ŵ2���h�I$���Ŷ^��<�@V�'������~	P����ĽÏ Ђ�YB�|SQa9���y��H_ݘq�]�˭�s�@;U�O����l0�;3��[�2�,�z��^�MA�����
���������<9̨�y��k�I����N�g�@� ʽ������t͜����YM�P��<$���'�-��r�2����������Aw&?ޠYHO:��Y.��$�2;���l��s!Hq�5�g~��y޹�҈ TM��glw�Bz[:;X���	��w2�w����G��� ��	#��d�z���VxQ�8��S��{ �l>D�4����ɘ�@����J(����j!��������X˹pR�8�ڡ����{����\H8d�Lk��������Q���{�Gm|�6�j����j�'s�?�H-�˱>'�tn/=4X &G�f�D�@�bPs���nd��)�z�R<�9�)�OF�4�l�x]��J�ֻ�M����C[.G�۝ܴiS�5�8�����$�w�`�V���F����d(TϠĽ���K)�S�#����z�v�V��UA����ΓB2�L���ǒ>�����olT�wTx4ϗ���ւ9��jz4b��ɯ��)u�\�.�C�v1�A/Xh�A���L����11h�g�ubn��QK#��dv����"�۱K�H1�����"�G�1�KA`Ŭ���)�2@A4�5��5��Ќ��@ϓ��"�#\�����?9H$��9��TL���T�G��Q�:^@�D�V�d6�����7�gG#"'k��":73d3:K�EY�3wee��K��0��z�b�Q�]����}��W�7q�S�2]tT0��o�o������A9>���%?~C���#c�f��.��O����o|/neF'Cqs�}nR�#�?y�^���U��5Vg�
hl�w+;��t2R��D�?Z�g���&�2H��j����~�ռ:'C~������ٳɓ�,�Y�����?bi9����쫫w�D��e?�����Ȋ��k����x{�с�O4O�}�����&�\n;:b��aV����c#/|��&<�J�iW�
��E��nX��w���Y�{�:�Ǣ��d��3���������K��?xE�+n�z˄���p]JJ�=<<�}���I��@t]�}�(�	ƧN]��J���i��h� �-����9Jۅ,��T�D��w-��z�!*y�.����⦠�Y�A���75x�|zGf�}U�*�$
�f�jf��r������b����ܮ;�Rrr��$"�x��
�ڸ��c	f΃3jķC�b��n��4�:�o�Ϋ�!�<z3�Ջ��Y�W�y|BdD�w\���FC+%MC��9����j�|H�c� �.�]���k���|�2�Eέ�p��c�<���OvBH�O�2�޳g=�F�\����ؽ2����D(�
/�<����J��c��LՕ��&0J���d /��vR�����p��^%�YJm�K9�7Q6~"��b硺�P��]�kq�y��� &�:��1���>�s���D���\mE��k�I�ׯ�̣aqz`K���Rg^�nȕ�pq��XkZ�P�3���u������������?G������Tw��7�������uu�Y��;NM �_o	Oo^�+c�ș���w�^%&8���I�`F�r�t�����?$"�M�1��䜌j��Mٶǟ��v?�QN�V���.��`�!9�� �F���0���p*�!��Xb0
�z��k���|3���r�4���%��&X��������b޶��|i�y����V����O��-��a���l��Ȇ�ߞ����k���r�i/�nc=����O��n칁���!�%�.|\b�؇ �BԲ�'RO�a#��6 �Yk띃R
րc����^��
��}w��2��+�SUU�zy�J&!�y�ڣ�"�
��23kGpY��a�d��Sύ�����c���|R��]��"����QVz�l�V]�¢!���J��FLl����9Q=�y<yּ�� �2a~�yZ`����ϋ��KV"�}��$�I������_�ĕZ���b�9w���Za�7�H^	�R{E�tp{�`_���*�����UG ?�?Ux���Z����S&4��=���n�dW���r1�ަ�D���Ŷ|��IK�ù+-�*���<���ٯ�	�]f�ԡ,���jq��/���n\����!�tw�q]�	��^?S�r�qŵj��'ͩ�<;u|�D)C��۽���==V��p�p�� ���v��>_֘����8���Խ�k����Qn���R3ۜ�FЙ~�\\M&6Դ�RJ��	v�ڠ��3��n ��Y����23��N�nT��Q,�{�r��u�^75�
�$���Sy�l����g���3��ź�����6��m�W�����W޻W�n�I;w����H 0�a�Zi��ګ>eJ���+�1��C��qv�6�u��R®�eS]������_�-�RR����ZB��{�>p[�p��Դ�Z뤑O�F���ovw����7w�O������F����ּ��QR��r�*�<+��bF����?.�Bއ�\�2�E6�Z�W�� {�̰ צM_U���Yp��(�>���x�;���}��8����y4�ת���fF
KI��z:��Vޝ�&\�-�;�� �k �Y��uF�����h
� V*�޲=^W�!�;ʶ��n��gP�KȜ���b��6�6qӼ�<�N=���x߷o���{n�_%-_�\xƻ���ZU(U��'3bg��Naam0�77��Z��	%�@������\~T����tpF����h��L�>q%`ډJX�ރ� O���9��&r�S��̕��/�&K�nnSp��T2�-���E���C��	�oj�_ݡKE�S�4��$J��o���uFa϶�;��+������7��,đ������aaa��*�uaPr+�� ��D/][��)Ҹ��.`��;�P�����i�F�̃�*Ο��X������Z�	�	޸�=� �]/!�fb�W�Ac�t7_$���-�)���tחv�:u��wX L�a���[՘�����ҵ;D�Z�P먗)?��[!Lv��B���}o޼I�OI����"]�!���,]���3k����5;�ZՈ�;R.�ps�l�H��.��� {�ݼ�eݦ�-<�uWH
Ϭ���[R�D)@L@����[��v���G�IQ��[h��(�����5	zX�EK5���s[��N@y�ETRQw,��|��x��3G���!� ��WP������1w��c7��w>�M������bM�$�NI�d7�m�8 �s>��f�z�f���l��,�x�s� �,�+�G�j��1�欨����{Sjq	��G�����ul����*Iǎ+��ٳd,&M�Rn������a6J���%���bn&�8V��˃��n�������&>������T�|�ҟMש��EM���C������p��)��~�����W�N�h�uq��#/�CN9��J-|Z����������jC��L�\��.�;U��fA�}ܪe�<�wz0@=&�m��_i�M�/<���7�c�Wx��2��r��7&6���
E7qqaKRO���^ęW��b׶V���m/��3��ZP�=(Le��� %>>��*�� {����]Ԯ楶�HFM�dnW�����Oy$��C2=M����>(�pǟ������0�a���N��9�����fW������J�����aJ��,5īg�O������@�8\�Cv ��_�b()?L�|����Z�g'��ĭ�Fu�U���xԸ���P�h,����x�;n���m͗�����g�/h���nQU�����>u���4c��1dV^d?�(��Ay�o�`Zj`�E�_��~
g�[A�QG��#jH��T�����B����� ���o����yl6��U���fN�Yy�h?�N0�ڒӷ],�q�(��[FJ�����"��(���� �L��L�Tc'F��WIdn��:W�uq�q�Ë��5����w \N0HE�\�n��0�1�۫�~�J��Q&n�t�,^m{S{5��Ü���{�;��kjl��<�V�1����Q�wkv�ð��ō� J�l�2Xw���@�^=C��J�I�����a�Z����$��
R�c���#�FT=\�[�}{�����-ʪV�q�?I�@G]5���xj?������߾}�7)l笛��|3�w9�d�v��Y�~����S�MR
i�s1S	��uӍ�ڑJ\�}�QX�Hr^Vt&!oª���x-
ΦM�p�G�{��~zLh�`l"`=��lT�0��[#mb#'X�!�R:X����0����I^�����l����qxL�e4��!����>u]f��*�|}�����l4�Â��f*��%��QG��my�qe1&-E�������4��X����S�۶G�D�Bc|ܽ����<�	�tn�_��i�-��.��%�F�"����(�(P�H��-`6��z�>�-X_k������6�5����mUR�}Ѿ��5���2�1�R�k����l_zwb��*S�l��n98E�:��[q�G�r���d�N�K�4?9]|	�+ڳ���#vv,.�
tX�2�]�_fK�`Z䱎b�mYU ��������q�t�Z5@
��YY	�yh��7~KV��7L!N���}}��̫���5��c�gx�/
:y�#����/w��t�L___ﹷk���y�8�j�D��4��eْ��?S�t��IL4�b�Q=�����V�޷D"�\��N~�4���^��v�8���K�峗4u� �m��4dѪ+�����w�G{C�i�KYhP=(���7	4?���:88�Վ�[��0D�}w�g�ͣsFAª�^k9w�K���Bb�n�����ag�b��|.��Lw��f��"����z$�,�H�"�e3L9�IjG�}g'i�|���%�rPJ���|%�"��֠sq�s� c�R���j�􆑈w�s(u%�FECϫ����x�ll�H>U�u�������X��6�ڵ�ť���&Ψ7���{�5���J�O �ߔ�3N�<��&7Qw-�cu�c�!�$66��A3J!`�������;�_LӃ�I��X�n��$n@�;X�C%�_	A�>�Jm�9z�M|.��bpHȝ
�i��KnL�?"��n�c\%{,�<�FL�������LK5�e�f��
��sއ�6�AKrӑ�=fݺ�=���qwD�Hn��nl��g�Z���*�␼%�v�wf�~.�T�G�$����ۍ��+ށp��<���*�1�I�EKY{$�׽Q;�ck�����L��@,x�b�NI��[� ����5;��R�O�I\%%�ϪE���;�6�ߘ��dC�S����Q�S����!	:\��+��4p�<8�3jYT\
Gɹc$��JA5�'�O9y��\���4����֮��W޿_�N7�:C�HH2���vP�eߍG#<�]:�I4����/Y{O��U|�YWE�c�!�:W%-	,��v4{_�m�HSG'lI����Z�~ʫo�Q)-XY;���,H��5��On�uy����6
��N\9§�6.:��{�ܰ=�z
��ql)��vG�U�o�ɦ<��1ו�ڸ7��]�
r�߱5����g��~�(���㚬U��^P��~��>��+ <������������T��[FF"w�>I}(]�_:|Ƣ`�D>�,9�&�7Q? �4Ϻ�f���V�$\%LbpW
E���Z��@ܬm��9�*�͛7_g���ҵ����sߔvԕ"l |�V�fi����W�j��������.|D��s5���,a�_�"�n�rh��PL};g�7���st�����[���Ԉ��'cVkd�o�4 �;|f���M�i������ ��"��<ǝ<АR�S���֗�xh�n�	�>���l"v֣�6�����[d����D��.5��̘�޹�����$��HUy��Q������3�q݃9O8��kr�)���b��U��gʰ� ��Lm�_wh=EQ���:��Oƾ"��-�r�x����Q
�J~�9�މ��w��REbvS��/���^7�Ng���1=s��H�e퉧BY�]�z..��J Շ<V��#��_�U�����	�:J��Zp%pO��D��΢f�#Ik���D��Q�(m��㦭`��ٙ�]_��i�h��@
�U.G)hXJA�IGqt��f�I��>t 8ؐ�%\�2�1'��g���j�A��S�|'|�P[6Q�h�Z��V/]s+؆�X)���BMH�t�b�Q��L�Q���t\�gE�z\L���r�9�[N��L�?4
?�c"~:�UC�i������ooԅ�#�]�w4�_�O�O�;��b��T=5-�:5�$Y"W��r�f���j�(��'}v�B��t���찟T�fG#*�Uf���Ӳ���L||BDǱF�B���P�$&�~Dn���$����P������	����7���|�F��h��c�F�D��c��NAl>]�Q7�%�D�ϯ?˘�ף�pk�|��i��]�嘒M�&�uE�Eužg�Y/��A���ě��bbb�r���}hJC5hV"���b��sP��L���*n��w�Ϗ�^H�d�<)8�S�.��/Ɉ�Ӏv���Y��,�Uz�챌ª �y���P����_�?TA��d�dqWe��1�^Gg�������¯�w����~'�qtbg��1;g�oGh���\?66�BB�A�<q�'T�m�C)�s3)%"��<F\�Zm��)�����c>WC�O|
<����]�����,����t-�;���|_txKl�~�v�?{	L�i���ƾ��_~�Vf���� B�[���?�����y(�@˱F'[�J�}I���x�А:�n�ho�n7�VB��������TtNWw�Ӓ��>[!9�YG+�O��D�2N7d13�Q-ز��ԟ���s&�&E9��|�й������W�ª��L�Ѻ���:T�&���V�z����:g�$���5n�+�n~����^Qי�F�ꘓJc�5��OEP���֯���!�+_������HJ`�+�B�r�써h�%��8�襜�o���~����Q�=.:���LN����F�)?��T�P�h\�sa�# �$Y�n3jKc�GV�͈��n|f�v��i��T�T<���!����Ց�%�dbk�;��C���b�˰����0>��L1��ЖFc�j�vߑ �W6*�f�=�o�8�Z�u���*:,�ڻ���Xbl��R�{}���,Z�(�?((����l����qb�_K
�,��A5��ss(lE��,�B~XV�Nq�����!�Nޯ�ޚ�1��UOff�����L;��3S�Ae���)�ha	�4�n4�BTՋ�ꌣml���"7R!j�_��S���M���<M;m���:�ݤ#��v��AO=�辨��u%۫��Yy%�#A���y��k����nX����M�3K�F
�t��K���%ܺ_YZ��WK�:�b`��� ��y��c���P�J�LB5?M��Y-ۅ\j�!�?~�u�'��8�2��Q�]�t�W��s���BSJI�[��77�>L%{���57h�z�zR����7:C�m�/������}wͶHb>�1[wk�o�B|�wW����v���k�Ν:rM�J\mD�7{%�����0������a�)��R?z����M\_otH��N>!"�Ο����MW�d{���>G-��FG��"�q*
�^^rf����gI�o:XГ�[_Df��UmkPҨ�;qTG�c(�:�k���K������S�X���
�݋�!~�e �2ԝ��s�Ƒ�M�SG&Z���Z��%�g)�DƩp IΥ�@8�i{P���^��f#L=�:�R����W�Vw���pt�r�퇋bߴ&���8�s.9$y�N�ڵk__K�]����D���!ž7��F-^�;��z��E�X,) ����8��S阘9_��}2s��۾� T.M;kl������Q����7�h���KZ=.?�q�ϭ-C�:݃�{�4�!�d�g'.�I��Z׏�\���MzA�o����޵%�+K�A^��'Զ6�6<�8��u*��5�Q���OXqf�sDa:�1e��`����WF(�\����è=�������f>�4#3�y�:J��7O(Q?�x�2u�+�W��*�qUJN��~������Y���H�[R^��V�[��k�����@K�$q ���9K*0��:!���摒�r̎e�c�jqۓ��-�ܞ��r2��֮����N�e:�گ}�(��ǜ���Ҡ��M{Hh�ɾ8�l��WD:��.�j�Zb�H���(P�4cX:u�3����녜{����M9�����k�E	��ϟ^�����3!�a��({h��A0����ؑ�a/��k�b$<<|����(pzvx۠3kk��g^�2����?��tO�Մ�}P�\�r%|�M��SeR�Be�(���6߹���6Rާ�yVd,��p!�Cr�e�SS��G�^{�J>E�Ѯ0���N�ϲ<�a�Ϭ���
�T)�_[0^ w���*��=�*��:�x�#B�VG�V��g;Kp�<�;� Gm���h��k>�;Y=b���й�ZG���%��6�����?+T��<y1��'Ȥ��*��RH!,�����K�B�*:��u���6q�_��۩��|4�e[o\w������|J�Q�O�c�\l*�.	���B(<���An0-��Y2�@�~�Ź�vΎ���F��?���-+Bcj��������M�V����TQ����ME��(����7�~��]՛�w˹�cT�K'� ��ի��2�V�O [�˄�+��ߜ�o;pM����WF;����A$����ڃ/�|�P���\L��L�	yN�m<��S�'�e#P�����V�Ѥ.^W�9���㧰6��V��Jg�� ��ʧ�M#�7�����������mɱ��G�u����������+.3f����G���j!�g��v�����\�n�'��~c�n����y���!:� �&(%%�^T�����$�b}�٢F�Z665�t� ��w4�D�����H>�ٳg�o���������K:�yl.�������zF}����O��":�~J�җcU�雖/_�'a	�]@���?��C9�J)��}0���9Ǜ�O��{�TXZ�f�k
{�m?�V��lv�� ��w���{��P����5m��K=!���y������Y��3�:����R��󨓴~Fd��an��{Ҝ5�N���$�7>���������X#�����]KEݚJ b�=�r�SnvH�vӜo��Ȣn�SÇd���Ә�Zß�&ݮ�g�db�2��� ϳ��:�@��R��y�&ř�(�9#�zO�2ݜ����ݜ�(ތXG�}�rS��a+��*�����Cz[�=f��V�	�Jڳ�~�YA¥]��VV���w��5���J�Z��xg�Q|�i��T���H���턽�aR�T�����7OeDV><E�6�}���S(�`�2τS�@�mE�ij�3��a�|�:$ں#�)`���q.�n
�ڻ�c#�4d=��7BC�5��xWϚeBt�2�vj�T��ʽ��s�.6G�U)�3�Q ��b"v��Ň�G�:='�Ջ����%�	��M�Q�s��B�OW�~�Z橣��� u+I;
���X��V��>%o�;��ڒv��L���.6�P(D�ӧ{;�'�������GG�X�W��>��;9z��� �7���gǌ�v\9��K�LL����+H�i��o�QJ�kYv�;��iO�w�'��A� oI�ۗ3n��e����:7Z(:D�Ŭ��W޳g}��c �Ҍpt��@���3ڐ���s|�,�:ِ��/7�����W
�}��E	?�,�C�bBw/H�� ˺�J�G�^!�z/�Txz�F<����#]`ް���0�Y�d��$iiiGB)RqH�nx�^�Jr��<��gΞ�@͊����
ɟ�/���w,9;��ҧk�l��;w�urr��ۈ�3��dq���g������uUp6Y�|ty�R�����gf�<5?(��ky6�����uhֿ��^QQa	�s��0����H���9�"�b����%ps���Cg�}G�@!����0<���lgϟ�7L/�)+/?؆����L�uD�
r�p���>���^()l���F��d
��<�7�~�X��y��|��yk����\HO!�u򎍍���u:VLL���J�J$n=5�}��Av-�ꮸ9����и�nF����5��������.쨾����TAv�T�4���W�o�w��.5�j��s���~%i݂$�� �΂Q��p���0$�PSG�^g�!��$���pmoEZK���.�g�m��m�6fm�Bz��7>�~��Q���@�% ��_�=����[N�����2^�V�v��SUU��<���A�)Z7�B�V�@�̶|Y��#��T)�6é	��� �)Aļ��^����(�ηm[0�N�_B��̘Vz��o������Ԃ�W�k%~�GL��@��H��a����������`DRRR�YFEy�?�	.ɗ�փ�������jN�(��˗R��on��-�YV�A���ו{N�zI���yѬ���ԡ˂:\��u������B�qTҟ�.����Q1�Qp��H4U1�`brGZPm긁YܔơCg���T���� �I��_6oJc�)!�kV'�6^�E��#��6�+��&�_�(� _B�\Zn�� �(�`���}j�K�G���U��*b����:��>8���sq��M���@���uJ��t���c,~�С�y����*2��-��{���w�NK�BI����l���p��BQ�xO&a����%#����;�v7w��%u�%�YZ�ݸ��&��M+�Z^^~�Q��R�t��[�Q�n~�P�~�p9���P�=�1�"�sxP�ߢ��m�j1̮���̶\YΝ�z-�:&1��XL� �{�\\9���S�~y[�(5pi熩8��&���44��� fjV16���A�,��?��a��<<!_�|I�h���b0�A�����kj�w�}ā���}�l'�b�`��Ԝ�qn�vC]� �9@�9c�-�gp�߹y��%�zzڧ� ���VЙ_��읰+��ۏ�m?6���B�@)��(Y�بӏZ����%^XA�_H�v���۽��V'�W�Ӆ���&��^Fٹ
eeeG��T)�RZFٴj��ү��B/� ��UN&q��A:�-��B]�1>�t�/,]Z�c���i�
][���+�Q�,,g�n�Sn��d���t^���W���#�2i�7R3G��=R����/`�EaeS��di+R��Ϛb9�w��4p^6��P���r�C�h݋��J��2���&ͧ)~Xͅ�@�<2=vb^����`��v:9pbn���&-0�LS�n�߿� E�Bw�];i�R��}�d��cSN���s�^}%Fl�6��4�Loȧ���8
�d�w~?l{a�L<��y�ȭ )i�r��~}�4�A��+{>En�$�8Hy��uZ�⯒9%@3��.5�Ш��f�+��B�'��E�Y��T��+���ʒ���}��;hSΨv����r�ԫ��; 2��9��:��F�M�]K$9ڦ�͗Q���+�^��+�
� ��A��4i,mk�����;_!����2���0d���Т��`C>W4xߪ����}'M��C��p<����Q]�5�c�`yB�[��q쿖gDWn^]�w��(?��n����0B��<���!�cU5z��d��ˠ�j�U���y
�י����y\o�pD&��,�U�F�ϦG4�>�Zp��Џ?n޲�}ѝ���W1F����B�������r���$�j3�@+ێ���\4����y,m����ķ.���{TYL.˼
0�¢G�_np-����������w�jYAB�F_��� �_AK���!�CV�����;��v��2�A����p��mXOs�U�N�ظ0��Y�D�D�߅/�)�9�P2�����Ɔ^�z5McQ�{��]B�� �XX���C���y�`(HWv9�'6/:����#�1����"���ѡB�[n?��K������p�e����t6��|����Lm�t�A��v��ST:�4B�翔������/9ܞ����b�RÜ,���ѿ���t9��᷻G,�n��'�.K?��jҹ�8.�xu��~�yA���vs.��+My<�B.�7�N�z���v���Ͳ��Kt�C;�i����sj���U�Qbtg�t:���j��)��Vq�KD�]�]:OD�nĴy����5=eb�?zb�◜�c�G�T士�=���k%֞ke<_���$���"���.�������.��2�~1ap�e���'Ht]Ѭҿ�O1����P�)f���EzZ�T�����T��������8�U�
Lmd/V?E�K�@b�����	f\�0���r�JX��ѯ!�:�j���0��.�q�2�~F�=0#&����0÷	�X.����U�3�3,2�q�u�=��x���K� ��W�nlg���3
3*1.2��3�ѳ'S���f���k�Z(r�"1�ta ���|UV�v)��%��s�>�*�,���\��bA�(��ۆf\v�\/,��e�}/��9c�b���_5��j!��Sn�C�V���2z-i�=�/���z�g��u�/+�}K�r���V��8��7]����g�/<cgx���]�'��`�f^7����b否�0s���˚ˊg�69#�����b�/���Z{��Jѿ��R1S貢�]-\&�m]K*�`<m���`��,aM�r/�O�?/x��ӿ|����-�l}h1Z.�ni�S���W��n�7�d�p�%}B9	K�cg���3Vxvօـa\?�D}�癋2�0kf�aMa�x�]V̔�k��6w�Ҿ���K���.֡t�en�Z���I�h��&�� $?���<�ѵm��|�6ʠ�R���-m~/���IK�.���3�g}ց���ZE�����=�o[,]ћ��܋|������_�����K�m�T,s]����L�C����t��r5]�G�;���q<�q�;`�^p�l�������f�J-�Qۇ.������Ӆ_�yI���K��[��k��,� y,w�J2�)�R��M*�/��`�.;�K|1��sY�,���=2�l�Z�'�Le�`B*L(��>a��sS��3t}�A���g;��΃���m�����4(��tY\ALcc�g�703��d�}�Ś�,,,����� ������PUT��?�����P�\��1�|����O�09�����.����g5V��d�i�Z�OB��-����-����-����-����W,ɲ��Y�����z�O��w��{�1��~�
�ʖo�?f#���[�o�����Z��S���� ��������-����-����?�#&�+�F��+����´�X��Z&��/x.5�?��V!��q'�c+��Ά�o�11[,Y���
�n*�h,T	��{$|��U���ޱ��z��|�.ےDl��?���rN&��ҘJ��l��D.��6+��	j�В$/��sd�%��7��23��;�"�c
���ma1+�w���q,/Y)�2��\ϸ����1nc�
F�\�_���"��-��E䕀'�Le�����L��-�ҋG߉��e�ϑ����������Ϗ=����XǓl�_��D؊������"��-��h�{�/�x�[���̲BEWWל{��at�97�Ѱ��H�ɯA�����~~O͐xt�c���<g�g�nnv'��B�ց��::�R������^_��ᝣl��{6�+�̵���T,�pW,��'��u��*��c9�(��0Lev/Y[�lV�"�saz�~hc�� k�4�5L��jd���0��d-
c��=6�6�+���y;��n͊��_O͞�������{{^����,ӫ�5�x��;�u�Yg��;���K����-+'�J�R�!!!'�1|�@o��[JpX�rrȩ��������MJy�݄��Y�ߍ����!��������q�0>_�w%n=�Xq	�Y�p�\l(��]3�D��JN�n�5/�OOK{dZ�1�7���#?ÃJvdTZ�Bں�A1�Y�7�v��K�FW��}���������Ƨm>�D��k�{`�ɮ���"n�Z�QeFZ����]j����ڰI���8g����I=pܽ�ݝ<�lp�h$�l�/՝�zIN����*����F*�>�aɼZM��V����y�!T��,WN���oq��da{�����5.�俬�ɞ�a.��"�O�(��(x�x��M��ZP�������>����Y�_�o���-j�C���2�����ﳖ$�Ą�c�]�,mqg]]�x�0'��_���%arx_�]>��Ŝ�Q�7V�jht���h����Um�3NC�� 	�LU��_��^�i������X�e��LL�����0�h���Di�,���.|���3���ljb����N���𣲈IH$=�Kj4�j3.�Ū����a�g�0���t�L9�kI���N]!��j[è�9W�#��1������Z]�/o۫�g�3�����,YZ5�̞�8sé��~f�1ƺ��Ə���<����B��v`zr���uC>�v�%����FJ��vf`X��]�1�[����{��^
�1��ˌ+.�\���e�aO��"ɐ%J�±�L��
�>A����]���;��/�EEE��J �VHBT)"VzQA@���  M��@("  MB�TM�$A����>�+���;�ޛ�3�{����g��Z�U��>��c�,lf�ど�{�q8WN�F����פ��Q���5�!qK:<��Q��>df��S{����n}�s|Q,<hN���\|ζ��5�ϊ�6y�H��n��C�̌��I����!�D��O�ڼNs���u��|qN1}T� Z8~�ڀ�ps�d_�E�}ƭ�9�L�(MAt?�m������OK���R��̮;�#�x���X5f\�9�b�v���u�r��h/�Hu"�v�`���۟�eqK;_��Ґ�	�+~�U�
5��z����Uz�-;eh�	***3�l2q'fW�"Z��\W�{�e �d�&Ց�C�544��h�;��dK�^����a������#���l������X�?���Q{�4ొ۷l�-��&�j\��D�hFn�WNf��؋W�I%Kv a��Y5e�++ǚ����^n�������ʀ�p$��r��ax�H*�����6�$����𙛛;..~m����c�����&��1�b �b��aaa�Q���щ�0'�e�#����
��V�=���S��ƅ.�8��H��2Z��PiJ�fQ`x��YjJ��!�����.��uh�Z��f:�wB_��)�c����,�.-̨��8�wnrӯ� Wjcc�\'��'I�	`R�J�:L�o����G�c;���ׯ��6ˉC��;���Ϟ9��|���lh�)�0��Z�;up�ɭ[��yV��ENM�0��{v�ݽ}[��=.-�c�	��Tmee%�N�����Ǭ�v�[q�4��l�ʝ��i�6��R�]�Y�[лG�"��J��fY��I
y2����!�ڵ��P�c�Q�h ��*�M"�n��&�� %���q�����M4����Q'��jMl�$7n���?ݒ�s3Y?:��:S!|&��\&����\]�Ki"���G�>~Tl�2�����엶]9FtĬ���F2�및�,�A���c�qPK���� |��%�fP����Sf���zNHC�M,Ź;1娇g,j��@h؏&�ӻ,��\�[��S�A�� ,S�>p-�6'��DI>w*�i�6� z��b�Z+�=?�NEQ@8 '<G@~�l�!}͹K�$��J�����]�(�����pK�6¾���\g����/1���Du8�#`X�]b �,�
lF;����6�Nc��ܯ�>�_*�A&A���p4���{@3���<C�kNP��>�mH�Ѣ�/�K�ǆפP�rm��6�XYY~���??�r~�UF;�f��3�ʦ��	�-<C�e�U2�kenJ������)����)�<
<�sD�a���fԮ ���������c� ,�ꕑ��q���ss��0]��� �/�45JV�g@J�Yc�v��ӫ�R8�3��ƻ���pE�~!ʠ���~(�{2�Z�*̥�NV����1l���M��)��]�r࢝Z��R��N&���q_sw��S��7o.Q:6�6�Ji7X)퐡����'�切�4�S�)�@OHH�B$j�GF�v��/@n��"��ju�.��%���@8ӥc�D���;��U��<�z��8"����L-,ِ�y6��g`of*[��|�� ė����Z������GK�����d�}ޤ�"ڊ`c���J���GK��^�n����aO���Q��ٚ� ~��nC�P���:��q���U��=h����&'l .7��&���L��K,��a0A#A�v�Omg�'A�qUʛ�)'k�F�� ��{���E��p�)E�"CK��&�P����*lԤ�~�2���@�Sz��Q�k�;�U�@K�j�8VG΃��r��s���E0r�v`��7O���\��ꚲ�di7�?Pʁ��`���O�*\6�*����e2�x�c&
��Y� ����*����L�1�iH@�S:_��:Ps�$+8j�����J��穧��8�l����M�Y>�2Y�p�ٹp���#��-:�@E����wg��~E����#a��m/n����O/�x��9Y�ʳb_le�Ϥ,�u���;\�x��ozU�[���������7���}+��̘����@��TuW�;\EUu���kRz�|��kN�q���F�|t�;�?Z��Y'
�/r1=3�mc�4<�S5U-މ�-Y��\�lP�N/i��#,,|�J�۷k7�f?5$��%�.���/N�O���F[@5$�����#��]��������::i�\�����:��` ��Z���/E�L�H}=�(�����.+H����)��9��~^�y���R�J�爍oi�U��;Oꤼc~V/�z������-6��z��i6��[�̞���:$O�J�ԣ#����0 �+D�ΡP��!)�uDb�X�Ɂ�س���M�ɫ�Z�����9kamt�%�n�_w\we-��g��W�k�x^nƍ��/g���Z�oU��^���Z��]�С~Z���}l��^��̅+ʭ*� J�QTvRP	~���m�~8�=[FQ(�T�S�f����R��ii�7�&�;�ٮ�\w��=���p�	�q΅�����6�gm��/7��eAh}��0���g*�F��eh�D9�AC[�.f�q����X�^�����g��<Zj.`Fげ��.�8��:G�a,f>�������%t���(e$��^��_:/o��T󯫻\��qK9].((��()l��Ɗ;F+g���,��	fH�'!���oR�����	Q���`8�+�v�3�C���l�[�({�����R��m�C�HZ�ڮW/żN:�-���� ��Ҋ�cO�x�GGF�޽� ..��/tUQQ1"GI��_�nw	')��n��CE��w4<��Ś���d��6DM�����4M��qo?�Ab}����"nd��#�n�sFR���QR��i�-r�-�ho�]���3�V\���SA3�9f\�n��ɏ���LMB��v�]�v�.�k��9}�n:�]5r3���N��^���I���������c�^�f
@u�4�l��G��_��Ĝ�%����]jg�G��'���\����YŒ#��:�'�9��B�vx���T���be�9R��ho���B+C;?ڛ
�ĳ�z����[ho^�NZe��+�]?��<�ia�Ww�-�u�&��o.�Fd 恜>�˙�b���p��̼�1��a\�������6������\`X!@����?���ڽ������mQߞ�b����<G�;=P��7k��,���h���"?�����~���CL0wYr6Y �6��w#�`��D?�!���m��oۢ�u��7q���������jjn���ၽ:��F�.]�����m�;[j��CM�{]�z�QZ�Z>G�5���#x�a�mz
�t�,�,�F]�gF·�I�݃��(���&V�&.� �-�������j�mx������g�ڈ��SSS9�T���4�;���[^�	���Hr	,]	�6A3�/�5���۲礧�6}�r�`M%*�lOy��>���F�[X�8��-��1��"UUU����)v,_���|g��t����"����eM������JB �	j��k2��FK��a2 ���)3+ĸ�8��	_�R̊ۄ����l+�1pp�:{`ic��ֶ3�l�:8��޺��@p"=Pu(P�@6��},�H̷M7Ebs�~�Yy+���* �?�~�������A�JZ�����@�Z�y{r@@ P�V�0�{�?+t����-Е+W����
41Lvn����# Ъ�m�e��60���w���i###mi��a8h	���p��b�:�]�5aC�R��E��Î�� lF���@�.7S�^�n��������$��U��w�`�4���8bz��Z�y�1W�R;���g�-�9�� H���IT'W������S�uc����q�!�������"�3�pX�<
l��9��d���\)M��
�&-5y�5��ɏ����R��>�!�T���X�X�?�w;Z↾��#��P���<�;�����k�.�V�G��2x���7�����H^��F{��J0�܇T�\�s,�̎Kq��3�6�~�FFR�5H��@�LWW+�����\����[{�\м9Ͻ9�s�*@�}wPՉ�J:K���"9X�:5=��f�L&D��v��e:��)Q�O�:ů�>�	��%�K���/�_¿�	���L8_|@��Y�����K#\��Yz[�<ǽ,��?�����O�=b��s�{{�^����C������=�8�pr�{�շYR�e�^�8�SMF��i��6�l��{eA5��<iA�T�e���>x�s�Hy��㿃��z~s-Yi	�Yvx��&�j���!��m�O׹�I'C�����hF�ű���7�l��8m׻(Iǟ�%�M��c�u����s��3��^�+�j���w��v.O��|^Y(��X�t��,U�	�(ɹ����^?����ɁzlGj�+in���~)6��[����H@��v�	J�Z�ꌢ�/�"��%*�n1}Lϋ߮$j>	@m�\BV�%-a��V"�,�����qn6�8�!��G�fZ�h�%��}F�8���/To��By�!Ӌ	OJ�+�7�<�8�N/D�m�#���;]:��+�Ul��*���Yp�Q��;��SW�1�q�-Z��(RaǪ-\'ܖg�d��w�N�m���Lō���L6���p�Ί�Pu��Jq�\�p�E��w��D�-M@���j�u[Y�7����d�Q �Yj�i�~.,����]s�l9�~��dȠ����oP�4�f�'�f����������\�B���n�4 X����uW]����>��[ˇ߸)
���U��\��V��)>Jp��IoN���s�n��߄%>�X"9!(��MKU�Z��sB�N{��d��Z�B2���I�)�nuu�8��B�Kv�${�	I�e���(�7�wO�5��b"�%'Q]�h��w�����Y٘"ϑ9:�����ֽ�K�\.��c�Itpc�J��般𳆲ҥ�?��(Κ#K���pF������ |��3*�>CG�O.��9���"Y���E(j�f�3�~t��������(}�=Q�4��t4����!�8���g�;|ź[����8{��t�E�sf�����}�����P
g�Gm�������<�ʂ��X�	-�Di���[kRh���udK�Dѣ�p��
���Q�സ���At�\@I��7nb\e�\kM6-������f�mԤB��Hw#:B��Ɉ�&+����+sN�C<�h&6R�$�ၾ����orD�LX�u���1t$�	g}��t�k*Qfi�f$�����4�_^���Gut����}�x��s�'�w^��j�t���\��̓Ϋ�%+�΃t�v8�^�Z��[j�r�����~#/'��,
J���N��!�����/t$EI���q;�<��[����H>�����/Y�<+�U>>��~i���+�TL��X�����d�9��Ɔ����$n��G���L8�dHr�M�;�l��b.����P��7Gad6�TJ�?���Q�����c._(�PB��3Ƣ�ua�a���kD�1(��'��z�����l�]\�4�5���;���#�#//_��T`��aNd�Hʙ#n�e��c����OʦϾ�r��	���]�,{��� �J���')�
���s� ӻ��_7�n|*DV*۳?����]�k��+�&�! rM���$��@�W���Rh�O�݉?��
x5z�қ��(�`Ei����?&���T�P�D!�rđ����N�{��4���ch��<Ԁ����*U�珡� ���&Et�"�D0+��#Az�ط��%pA���)�?��]*�#����Y�}t�t��協B����A���o�AR�Q:M`�鞣\��y9�.W�ߖK$/�_����Qw��yxD���c��s���Ӕl�e�,R��	Q��- i���&���6�Ku]�7���4y�$_J�dw�B2�H{`(���G֓ ��K)tȪh��8���H����8#��� lXȅ�%�6�7���o#�WG@W��m�gu�mAJ��XVG��QQ��:�(���l����Y�G[HP���y���,8{OJ��H�6�2S�ML�K���^ʵ�OAk�I��갤��m0�
}�E2ӐM��SK��E!�H^�(��f�}�j�P|Q?��{y��]*��j���&�4�!x�/�E�w�%�"�
��.���U��h��l���P�-2<���$�oNUK�_T-1���Ѳ"��%V�/%r.�d�<@���ƽ�	�IX"5I+����5r���x�6BVU�	��\�I�&	P&�:v���H�yJBV�n��Ra�:~U�f\�o���k����!�=$��-�}A���/<��R -�Ց @C9B|�:��^��z�����*�_;0��mp�*U��Uu��q&�ʺ���KG���N��j��R�lR@ ���A4�4(2��� :��¯ݧY 	Q�]*�)��?
#�XJ}>�z��Y@�	�]Pu�o �=��ʯ �eZ��dQ<w�y�n`����A�k���	�hy��d��Ҩ[�����J��y�h�As)��L�$aClHT��~ع�'^j���*�]9�@謤�q�z�:�<T�S���3��~�IG�%�Y�6��{8l�U&��lC���:�fJ���)W�ZGg,���U�>�[��~K���yZ[	y����xD�/'�$����9��p�b3�_o�6<���u����Y"�B��
�~��Bc��
�"Z�!4����3~r���ʐ�����c����^Ū�tV�9׬?"�at��� ӧ�jgٷ#3\�s�J�nX�,��f�K���(���4��p*
�j�ي 9NMB3�ٛ�=��ܮ ��SU��{W�2����%�9䁒t8%�'N��[�_?Ȟ�%bx��/J�P1z��< Uxm�Z�����X���_LdE�Ʃ�n~V};/�nO��{ �5���B���r	'�,%��k���8Tr���pe�i�󼒓�5*l�K�<�3kG!ϙ��,��N���9gn[�*�\����u?8�+��H��L쓔S��sj�#��i��Pf�y�d����uh��҆[��D���Uc{=G.�y������Lv4�^p���_���-�Od��.�T����6��s��a��{ف������vڑ*��^�e�ʠ�Θ�up���hR��b��U=Duc�o�񈭼6���[��ߤ�R�o���t���W���+���b;7P#�,�j�ky���A�/j-i�_n�5������`���ʎ���	w~�,����[;&�O�ͭ�h	��7������F�m���\��dgΑϥ#ƞ�$[n����]�'�ʐ��%b&���|�"1[�1�ve��o��n�dL�V���������<���n�"�/���Λ��ya��q��r�)�R:Bl'Pz��=���w�]�2U%��g)�{tZ�͓:l���nO\���a�Ϸ���{A�r�#�� ���V1�`�UЌ&J��A
�˕+&�mv-,I��[��nܾ��;�Sa����(9���dU�G8���pl�E���$�����{����Y_.f4" %r��O�� �C����}�;��F���s6�C�Y�'���Tl�p+�I�����1�����g3u��"z��Ny���i�%��|�.�Ew���h	�L�M�|6������~�׌&�|C!���?�W>��C曟��U��5[�S�x�5gS� �FDȦ��BE�S�&0�%��=D�ﾞf����C�I�"��;J���;�DTU�X������3�=��:�����=GdU6�w�x�N����9wV�o�y�4i*5���b���Q}�E��܌��
]�t�@���UĿ�o�- d��4O��g�#U�>��|�v1۩I�V`���������*��>ݢ�.#Z���/���@�꿚�]��� ��Nnf��>�d�q
~ ��_�J��s<b"���z�J�7	��P�Oأ��:uχ�y(h3���n�og��p�=�����Ǌ	�4�-��)�jfʟ)��+�
��7�lô���c�_}�^��g2�7��d{�گ^���j�3�����g��(�_9�%�-q|�JPM*���8�戝%k����~�%�4 �$0� },��h��Y�şOK�;�H��N���m��eXs1E�*��>`29P7[)^�~z�b�p"W�&�	�i�`�7� cw �l{vL<,D���w��'�'�o�����@hېjc�@��F�ʥv���M���ǘ�Eop��lc�,9EKܠ�a��?�5OM�J��Tj��{�vU`IX�{�i�L+ã@<�+
6�.�8	Vd\�i��ԥ��h˺�o#2�2�K(l����	���,ˠf��,g��^�����R�����T.Z��G�����p�sߧw�ݡ�|t��
C.57L�Q�߇�9���#��D�_[�n��	1o�e\�/s˸�� ��23��	l��F�b�Ri���k�e>���j����6?��C�>�����_¿�	��%�K���/�_���	�7Q���Ф
��x���Y��Ǔr�ْc1�n+�SlkD�����e���7٫s���I�����jM�_�}D#�?:KNiJ��x��qv��h�����țO������a���,���_2���m:" ���%�Z1M�;�"�͇���F�D3�Y_��3ȦӁ���gi��Mu�`��E�U��hh*��ԁ���bܦ�H�/pb0|�T��dջמ\ng��Ùsݽ��������Pl�(V��v���u��}�6y��0ف�a�ӯ�r�>���R��$���^���XN �28 N~�8�C�/��T�k��Q *�(�5�Z��BHc���P��u@������͖��^�`�V �%�� H3�=�۷���[u�����A+����-v���|����/�ȭIx���0C�+�x���uz�������:�c@�Va�Hs}��74��!�>q �J&�V�V�+��o\���>�"�Q���7��"��5Qb���
��]�k�S-�$�����d��Z�k��;����1`�e������.�W��c�Z�ti �Y�5��"@,�m�����Za����jʕ�}T�! 7��P�%544��&�B	���:i\$ o_�k`��g���s��uՐ�V4z��ݙ5�F�uK���u���� 8�ϭ�m� k�����˿`��x��������5$P(ּM�}`�u�4V�~@ɿgMF^/ M	���}�ݏ�E��r�\g��,\����\f�0`"�.� dJ��7��c#TL�UR������%;
��=�{���D�2 ��)v<F�q �lYwp�E0���j]�g�3Q�X���g�>N>[�*@��G�$�{��ׯ7$$%���;�U[���l���7@�ZO�z? 8eBh��u��\Z@.n�5���D4�5�C�Wa�O�ɒ`�HE#���T$+ p� �+��q��p,Z�5ܫ6Nu10%4k\M	]ӛJl=�. ��C{�=���CO?Y��X� ���]��P��`x��G�D ��-�i�ϭ�� $ǁ�w�7P�gL���"O�C.�,4;�Q]�|��a^g���*�w�z3qîgJB���0F�Qk�J�}��N�H���o��?���د!=(t騴J�a���-�%�K��lE"��}N��a|��qMg��P|\���Z��ޑМ��[;"nd�3���M�����O�������s�Q��B��
��Q<���Rɿ�2���/ÿ��1��?B�^�ߘgH@/ؒ����[k{;V�<� U����z?��H��v�LNMM�,#2�h�U^��7b��ƙʐ����_�0,������ʲtrBb�@�-��xxj�� ���@�n^I	OKK˪C�=����� ��~�3)�,T��_\��?I߿�3���
v�JJJ���佪�-##���d��R'��!7*:����������Ia�M�R�(�K�)=H�����f��5�~�&��K>�]hl��֒D�˂�4=��3EhA|��`û�������;�s3$����,*<'����D��2����3��h�TUU��XsMEE./�T���b�����-�,��O�>YZY�T��8���եŢ{6�|�<[#���ttt��x�����~��4�-�<�����0���/��ug#�PO&_��_I�I.0r��r������X��veFt�ѣ�g��#���ܘ/��%��\U�xv��	��u�s��7vw^~�q��89�&�%�l���o;e�U5�97�=?D�HNLI[XyK�.�ƽ{p��zW-,�B����#V���Θn+\����ēG��ƿZ.�-7�B��}k��6u��;Yc�
����I���gE�ܠ1p9��ƙʇr�3�wA�����Lk�Fcn��Y��=��;8hu[7h��A���Ǯ�x�<�PEA[z��ֆ�^rCl̽�$��,<�jh D �N�Q�u%%��ѱCYn�	/����
dC"_\?������F�������?��^H7%+�Xp:$e���{NS�c�	����̾�+�]����^3�p�����1'� �HL���
������;,zxtFIA�Gq+~r�"�p+�;W&	&��*4;�E����ݬ-����Zj��-n'l�}|p3�n��[�z�|:�Te���iv�	���0�Ӝ0�<)m"��#���gj�IT�*���ɉ����s�sN|��h�ąh
j��D&�"�+H�F|��&_�����sDr��g<�]v���IH(�{��"}w���qN��A���"�W\N⊷�0�nj�((xq�G`��������{ˎ��d�w-��x���m+]	ߓ��́�A\�$� '"h�a��LQg7�/���%i���!���j��xe����[��}��+έ,�um4�>)�d��m`�p�le�����J��d����L?'U#�D������\�D�V�{{�o/���*�:ݹ�t�cՇ���I�!$�?r�W�T��G*#�d]�ud}&.��#��ׇUf�!;�_%J�IAD��;L�W�C$0)�@���])q��&�+�BP��aC3����]�$�?m�+OGr�V�|(��y���_X��mq�KO>��5[� 7��[
��o�zJ{�׋�������J�a�U����nC���4�Oq���*6���.��Ы�H���~��I�I��*U�3�N��2����BE%�ӑA���~a�/�h�<�y+�����!pz��ܯ�/oٴ���g��qI�)q���3o��꼹�и����V�9�̅7�D�%�I�<1W �8L���f�nD�-��Uyɩwp�͏�\H;��������O�M�����_\bk{c�*f��՞7eU�]���7y����c�Q�u��x�
�w��q��ȍ]"%��VjJ�s���v+�Z��F��A�a �(��t���B�.23O�OU4==�g*���	(� 1@�Fn�ݘ��M���t��w��Ê���C��^��K��g��k�Vxz���5]fBZ�dB����ځ��f�����;�{>X)�^s�|}���m����?q?�ī]��㨅vHk�O��K��~����z�����,��Xlf�?É�)�]g����'a����3��֬޶���3�s8����R����Bσ�*_L(�AQ_E63�6�=}��
�R�ZjB�+�MRvGøQ;��+������M���qwk����v=ͭ��C{e�/%U�Tul��7g�i{K�m��6�a�����ܾO͉�.a���6W�[V�����{#`z���&

C�T�//%��a1��	#�Ǐ�#kTwF?��ִ+o;��~�w�_Sw��G�6�*�V��)��o�MvD��M���֎�D�L��>��ʻ��s��?.���w4fRմEm��I���i��������L��M��۔ǿ_+�n9$b��,¡Ӛ�\�DB��d��H[��r}bO��Xe8��Z��kl�Y�s~���ȩp(-���o�������<״s�B�Rxi��N/pȭO�;8[~H1Ǳ��j��T�i_i����~Z1�'���CH�ś��?@!1������%���_����5LY�=Ly�ț����[ށ��Z� @��
y�{Ə���F�Y%��w�:��z\�«���l�y�?��j��sw�9D�f	�l�c�8�/�R�++8DT�.�X�\��T�\N����Dɗ/UIi74X��l�/49)��t]�*���M�z�ۓ⎗�ؒ��>t������~O*"|��e���od��u`�؆<����G�q�oN�?���#��knS���`^<km__��).iף����E��<E����3!pc62��͏�q����JG�8��X��avN�ZEv�L�|:������@�1�{��B��`��F�]��u��_�r�����و�\z�ԝP��e*~�e�f�������⤠l��>W�ۙBkS�񽐔BIH���\�)Qc9���,�w��"�[g�� }5Oi��R3.�**����H��P}�|�L#v'�쯺��8��N�r9[�X}��۷���V�I��TK���A�P�T�I��&ܭ�f\7��첩�0{T4��HBJ���}�Ӥ�����Ge��~�b��~kʭX�j��� ����x�9�m!Ŕ�J N�N�d1N8* 2R>�v�#Mw�a穂���+� ���w.,88���D���je���w�.X-i�<�e17}�;����/��pnyQ�k�ȧ���8�ږQ�M
��Pp��%w�ƆO�]%�գU��b՞@�pq(��ߣ>�Q�]�6���n�L��jG��4u �`�Q�]=�j�dd��i�K��o����\�K�W���%6���iRR��9G'd�T�xyx���wy�pb��)�Zsb8��6������Q�p|!�jRR��6o��t��k����dk H�$�ʳ�R��W�7}�?����� q�c@���l<��5���T���֢î�n<E� QY�߷:,V�r�`�\N��W��4#����"Y�>�*,Ǽ|pwG�����#���^��a���V��]3�|�N��ַ��C{�4>�%X�p
�`O�|	ʗn��c�E�4*�o�i)���Ywk]�Uƪ�N�#[��+�٩i7�޾b���������M��|	�wU�6W�-�T+l&ʲ*�~��(E�2��U��P�h�̌�l+0�����N׽a�`���QI�m;T=�NZ!-Mˋ"�#?I��_w�-�64	�|���ۿ� ����HpJO>sI���Fuff�Y�A)���K��]�'��$f� a�x|�T^��ԉK�(Y,��װ�Xk�\~�p�6jD}���]�l�R�~tm׀�ٟ3!�h����b�bN��yt�����m���ح�=$d��x�����y�'$��%YX�w�+V0лyЖ-f{$'���*��h���;�~l�Н�,�a5���'�5�Z�]L�����/"��y�L�5�g'�jK��dv%*�UWx>��?� /��#Y'@K���YV/.����а�u<8܇}��_�΋7��c�_h��F����iE
��1�ͯN2�������a���I$`��}#[�nT&y����\�����s+3�z��_`�BО�?�b7���#���Ğ�N�㕕>`]@E�WMSA@��{r��r�~rk������m�So�ć3�D���8���U�r��J.^n4�~:��,����Ao�r���2 i��P��G*�&]$V#���q��IǏ& +d�אoJ�ӯ���T�"�g��Ñ�i�@�uhܳAoZ%
�`�)��'@g�Z�D��_��	�a|�D�]Kμ*�Qԝ��6�~0c�8�fƒm-���3B.>�;���y�wl;["g�SI�ma�-�6�-O�\��v��(�\	.�(de����Qs��{�Ev2���(<��<h��M���ٓ�L �&_VA@'ƍ��!�>�?0p� �R~�5۶�1RoL�#�w*#���z��_�B�#� �Hjm ���,�Rۯ�Z���0����c��>s$����)�׈�?��@�v4�,a5�}���#N�H�G��8���WV���u�6���������ؓ�_3��<�Kj��<'7��l�5[��`�q 7���c����&և�32TTG��nx�s҆�2�nN@`@�H2|�:�<>te�R��f�y�.?,p0�S4�\A�	v �n'+ې����"�vݹ�L:��.o�H2�����T�����j������Xr��-G@�CE�p�+���&���&�sj�}��r�:��{���h�N��.H��U�������Wc����S����D�����zc�R,ù�Vc?ը�;
f���P�}mT�rK�\�a��7�=�k�ݯ��eq��̶'����=��#�0�2�3�ם~���sp�z����$��t��.u���݃'R���^��0Tq�����L���go��ƶjhb��	n{Y����Ր��M�MON�h������綐����&�P� �x��lM�O!y������5׏ ��e�o�1�ĄKUώّP�U*Q��7�]�V��q	��r#�\�`g��-=ofb�y`�`�s��;����
Vb�iK�y��`���Ԧ�J�5�-����J\a�ڍu�C;(����~p��a�t!�����e9� �u��V�P�{��p��ǝ��-�1zH�|,׺��I['[��Ĝ�ga���ϔ xGĸ�0�/��z��n��!#7s��ԁЧ8;w���Jd!�F����1���|S��%���'�*�'�����۴�Mhb��DM��h�21+� ��������n~�.7P�l��0��S?����j�l��
�'2��Z���ees%Rs��[/��>M�ɱ� �}4�p�#g�ޯ�#�
�S9FZY�?mSӇ?�O�PE� �?-Es��Q�*cb �qV��6�L��m9���6�z=����&,Lhx�ơb�aJ�	8/�v�"���g��� 9�۩��f�w�%31��E�`3�9�wTLt'hU���݈��rb���.j��4����A9"�"���c+�7�k5$�ϑK�F��D�w��4+zi���ٚ�DZA�	�^���Ø�um�y�ʌD�늤�̙�Ǎ������d}#�W[
��ν�ly���9��1f�Ij�X&�����U�C?1|-I��"_�%���wZ�6�s��*����M���5�2p�q��K�T_�c�b���6{�Q�������)e�
/aU��[:3B�a[z�����򟐓#�a�%7��t�����(�Ă\!������JP.�景��g�}��NW�앓�޳���O�Y��@����$9������v�C��ގ����*S��/蛜#9�{���JU�R�i�_�%g�w�'��8�VAy�GG/�86L_?"��V:�����,s������O��M(���WU��@�B0��g��n�Q��eJ��J�B'��r{��A�'A��i��U��:�����Cy�Mn<�-'=M���ت�NqD���m���_*��|�!HҶ�Qe���l�2��Ⱦ/I�b[5�u��T��2hi���C���*:`��yd0�����rC��e��$e�/����8fr�U�.�E[r�m$R*	�RcW#�o'��ʥQ����������ۏMݔ�h>�r+�}uk�"G���d���T�Ѓ2[^��'%���Rה�D�����e7�b��^1dN�[�8m��g��t�SCN#��-����I���2I��Ҟ�'��Θ����v������d�ݓ�]�l��5z]�zfh/^bW�YP��6����ϵ�uuu_���1oG~�P��b�Q~y�v{}�����+jC6�*��F5>��Z�az��J战43j:�S;2�h���i``���2Y���͡s�f�S�h��ȥ��b���vX�H��|��4�ZּՐ��8S���/�Y�i���4�C�I]	��$�ݱEL��}��8���jm�2��d�}���O�ʱ1t�����xu��m,�D�L�@�p�^���8?�C	ų��+"/.+F�r}V���yc�)��UB?��6��>A����+ŋ�VR/��Y�6�W2�����ݡCw7y�>|�|C}�|�O�!����	/V��}�0�O�o/�K͜�-�Q{�7�/��A���9��ٹX����:v_F�<�ǡlw��z�x��]���+��) ���\ZU�t.�|af���\쳨\�Y��y�+��Ǚ�-�n������"���q<Kd����gJV��UWe�C�E� �e]�q����1��:yO�����n���_�q{d����)#�܂fH8�Ȭ�!��6��6Y�B�]�*�q��#j=�!�F��=�ޥ������ ��`7�S�(��CQQ�dׯ�����$�$�Tm�Ú�4=3�6a��lc�}��b`:�\�^ڧQ�ֺd��2S�u�ǝ<���+�Ki����:as�����7�,�+8jq}9�O{���z���l�f�c'��XtL���b�Y3k[���+3? �4�dc7���A�F��o;\xD�v�ӼABzj�G�5RUjnk+��v��UtWަ���v�#$>/�Z�~����OB*�����HY���ڼ���\nJJ
)���G/?����y�U��!�B�a��{�Us���A]�j�vX�;���ni����j��/�C1A"�ԥ��V��U����{������D˪���Դk?v�����7��Aǉ�����3�N�ǆ�VT�B*���2b�Τ������Ǯ}�"�X����`����{����%�0�bwU������w�G;�Pd�ڋ��J����c�(ΰ~t�f���Ž���7����_v������T8�ځ�}�;����.�<�0t���m��*�s����'ϴ�� 2RGE����ia�A�TP�O�?��~�an�T�m�K߱���6��cP��޾�PN���[��]Ʋ�$R#s��[U�{��t��[��n���^;z.����N���j���C�i&%%�l��r���܅Ґ"����wE�������'"�N���-,F�MϞ=��!}ثfmӿha
�8kH�ª�л�xƋ��_g�e��cc���F]���V\Wb�zX-'��5J��ٞ��������{!�ٽ�ϊ�s�pU��^�����=%�Z���+�H�/��H��M�����/,B��s<���l�}dr����|��VwQi�v冽vխ�gF:BO��Q��g��A\�?t�U(7�>A/o#	�վ�ٗ�=8�JY�s��~{޽�q��o�L���%s�G�Z�	^��K����i��r��P�$��i��ǆ؉��W����׌^@��"��1Ӎ�-3%<ۭ쎍RR�ÚY�@�����r1�&��+�J��RE�h`��G�=���U�.�?���W���%y �T�n���O�lWW]��]�'��W7����2��PZ7��\���C	�C�$���c$c��������y�a�������j�6RYY�1騅{���J��z������a�}��/�ɏ�l�N�)�V�t���W���ś[ޛ��D�*zꫯ@���.�/�d{\!��Ϸ�`�󥥘�AUꊽv�Ŋ�M������^��&�%bK��P"�]
�D��,--����J4�����|���\*ب(!�bI��i��܎��f��CR,z8�@���� <�r�.:�����d[Ntۥ1� gd4Y��|lT��ݏ��YN��5Ca�ͳ�� .7W<�x@b�t�U͌E�D����l5�<!�2�̻�˜�h���O+Y�w �жoO��J��r\w����=,{�}>E��[TJ;�C�9ن��~���ݞ�����f&٨��B6(;2���\.��9].x�Tp󷝡V:�)���1%2/.�Rb�A�l�˺=�ȼkęېd��w�xei�(�U��I\I�^��Yv]��5��bG\e��^)7F�����02�.>ƹ�o� �k'�Ge#.,,;��+�ɽ1���%�ȅܺ�;�����ש_���
z�HN.E(��h�p��N[(�fn�xV`s������f2q�6�c�F��x`��H���+�<�I�n�������nBG���;u6e�01!���P�T�Ʌ�K��l���h��=��֍,G�v*;�@�0q����`�Ѣ��!���DtB�m�w�6B��p/�����c���� ��WfyԤ�^��e�{�8Z�T;�_&�q5���?�}��j�����aQ�]�8��� (!"�#���R�)!�4!)(�!� �9��H�(1RC� ���y�������}x73��^k���=3N7��xPMR�7W�=8) �:��Z�8� N`��`��]��w��4���s^?��th��0���{�O9��ӊ"��Ĥ㮘��_�e��q���K��Z%�og������z&L��)1ҍ��FUV��K_��a���LUP���=�ሺL$�[�����z����/�y)G�(^�A�X}��NN?���!oS����4���d����Լw4U�J�����'}�
���Z
ԷM����Z���n���S)+����[LM8i��zq�ߚ�W`�ssM���MՉ�?,��|�9��)�A�b�iŽ�I�U���ƀP�ȼ�1>��!V���H|���$q���5�z�cL�	��c[�����fa��#+c����\駄�����&�Ɍ����!#+�^�	}��8�_vdۉb����!,]5/4T[�Y��N��D�g!5k���������ϣ��̏�ZP!rb�rX�$τ�s*�ӹ7s{>��kM!���Sa�m/�J9!���;�kHaJ(5�� ��`{�{���1�+��7+0����!ꮑMeW>QHH.l9��̘[�-E9Zk/�����b�W���o�-;�T.&[ ^��)i���(�������{�O%�Pm��" �'�r��j��l�6��AOGWP�-ގ���6����n�G�X*Q���D\�]�u��Ed�'�'���;���:�^���F�n���/�M�Z3B�9+�VN�x�V�U@�4�ʹ�AV��SEo՝N�@9*�p~B���39��������n�pF�k\�OM��_rtt:��\0UY�ܽZ�(|�j�V��}����iFQŽ�z+�%h�'��tȪ�=�11.�Hx�Y�����N�4tP��d��5���b���v��w�.�K�yF�����kP��{*�*�α�n�#q�]�����!�����C��XCz�v�\���v��GH�f�4e�ͻ�0�=��r��=�B�qwp�;��d����8�~�r�r�f�?O�h���c��#<����\��no;)**9!�����{�u��Tx[���巠�ǔ�؅Ƚ����{s�V؁��p��4�*��Qjfa�$�M�����T}�`mY�)
��E|#(�������퓗ܕ }K�4���� ���ƹ�r�Y�E.)b�7�꽂�������O'��^�?�T�5��iw�`n���ɠ\]��6�+�
���:��k�V09�����VA�0	����B��=�t��={���}����z��A�A�x3�8�=�����A�ttI�ɉ�#��h�ۿr52���F�ӄ�ZH(XV,�6O4�m��R�{��]=��dUyhSܰ g���ߣ�X��[��N��S���)�{�q�ـ�`�����1[����<5<�=ߣ�����9*+* �-襻�i`��=���R���q{��KTg0)�����£&��kO�<��-K!��?d|-���.����64*����=T�-ju�����ͷgT]c2}4��,�#\l�ԩ���/Eq�+�.�T�*6&?��"B�'<�|��/�a�i�!K��n]���T�߰G�c�O�d�J���L�4��H��\���j!(����D5�"�,[�t�_�j�"3�F��O)�e�o�̯U����v����qZ�ʗ6>��,�Uru�nS�d}�H�����c2�+
5�$�im������Rs��f�9̻�ʿY�Q�Ds�(Vk������b��H��i%�OȲT��[��iB��@U��NŊt���SM�`0��Z��Y����G;�{/SN2��O֬Z�%����D���m��j�DW+y.�������KXn�>=�~��8�{�ׯb]ïBz]7�ߑ�c5�,�{��5�[m4(Mo ��9��b���[�5�>�#(�j��}D3�S���3)�OlZ��~<=dY�ͽ�I�#�.C���C_]��y�"?�O'����`AK�6z�y�|�w
��^�k	�z�PV0�7��r�p?=��5+�nEI�$�g8��=�C�18I�/�M�ס�_~LgaEѿn"���Y�5�X@#Şk���va�����1@�AJ���C�Cc���x�u5���Z�S�qz�V���r>tR�� G�;���
�`��"�N����7 K�e��L�8k���Vٗ��u�KC_X�6{�K�e���X��s���!Tĥr������r����i� 	{�Z��U����Rd�(��QZ���X.z����c'='� އ���R���/|Ò>�����Jג+�|l��ï��)'�9��Z���x�k]�1�E�:@�� �`�J�S�72���@��X����>��gl*u�hg�w��-�}��4�Vt4�'�>������
����uN#������D醾���� �b}Å�b�����2OP�.������ݕۋ�}�{�Q�4u/q�f��Io"י��0P���툝�5U�S�5\EÎn?�x�H����:�0.R&�^Z��He��GT�L���F�E.���T^xV~ڈp���)nzzz��t%eH��[�����O�ڷ��h��W�����[�K����-Yn�(p��� �CK�&%���xQI��P���t@��9:-�D4��!B5t�F�t�l�~�8�EaC=�K�����g�M7PmUz�}|���A�Ɗ���Q/���s�V��y��sQ-���TXg Ƀ�,�!��c>��S�{�ز��b~�W�{�b��>��/���� ����Ɉ�������f�y@��Qn s�����>��_�Rmҏ�j����t�Bq��ɔ@,ͺ�;m4�����x*�$����L�`�RTo���V9�>�m-����9�>��ܝ�0�4J�7�X$$��)'/���~4��ü��p$����AS�oZ���w�e���?tW�}�֯t�	D).2� ]����C����-s�ĵ]�Q��*���N��j��V�̹Oj+�k��h��`p��9���+h�Ҩ���	O.��}��j.=�W�ii�����ޚ�%Уh(&� <cp�5c:�2n�� N�A�"��0Z�G�L���*��O辩H�mlSSI�,�V�x�Z���(
���z��Yo$I��KN���c���sF�k�	���|�&���氵ӕQ��>iz��݅M�FmU����nE,��W�����H�q|�i@�h��4k�8���u�o�U2�h�XYY�	A�`��g��~T�PD���4z
�?�=L�&$bA�GI����]�ܿ��^
Ʈ�AD�Zn.�8��c(���o|B�`4y��un�S�:��t�����T0s�j9>�X��,P#��y0�-?�8H��S7��S���^䞯;p�ݢs|Ş텃n�Z����Հ邏x����LB>�zy�?����V,�%D��V�G�dc<�d�AE��P�t���ISrr��ک�օ��v�������ܣp|t�h���A+��R�/:�N
��uP>2'D�]����,H�N�y�8�������XTX��"��\���j���l�9i�i�L�᫓vMi��d���
 4V��#��3�1��W�!~ݧr��5'���޸���Cxx��ۆ@ۯG���t��t��9�0�7�Bэ��|@�q'''��i�)s񣱸/_@�?�LFb���ht?^}�V)��p�j��_��+��c�N�-�x�)��/�S���^g��P.3�y�5k���R��2��^�%��B{ �4� %Y�=�*��o8Q���r�Թ[��(SN1(>��O�6Z�XZs�`��F�Ζ^շ��X�����	�%"�ܚ�7���� N�k?�5.��~���M�ŷ��<�T�����I���^�P�I��צ��v��nBmg
n��K5��1�X��Y
7���6utZg�M�9��5u����CZ�k�Y�@m��GWO�kuCθ��Ԇm}���2��{F#	@%������l6Z��������̣2��	�a�<�GC���w��vv����Ӷ�!K��)s�9l=T�m��p��p&2����9.����]������d�u ���ʮ���@b���=��+;��B�P1�Z����;�웃r��;����M+����4b}����^��.ÓW @;h�����5<�3���o�}����Z������\�o�ۻ-�4�� �u:r�tr�9Fܖz��	To�}1�V�S�%�_���<����b���
�C�U��c]V��}ҋ� D@�'z��Ժt�sh~�A_Oٗ"x]��2+�I$�X�]�ߓ�5�%*C��-TVh����������w�d�
�{u���Q	�$&X���4Q�JF�^K~ʆr�?>�?�������jBs�]�f� F�ـ�z�(� g/vwdo=k�l�L�S��.&��ATgx �(~�4ou��)�n~�;dI!��8Ȗ�E�(v�ݵ�e_��rl�@ӏy�G���Md~u�mO�]t�wEN-(��;EޞS�Շuǭ���B��� A���H_���JՆ,(�����'����@1
����ǚ���3G�����4�Q�} ��9q�M�X*���e
gsD���3���Ϗ��{�c],�y03�j��s:V�e��6s:��#�1P��R�S��`���BR��,U���uٞ�\ّ�I薟�����*�Uh�
�}���(������S����8�fh|��Xw&�<�w�x���=�}���x:��ϭ>�"��S��y���q�jV����c�}�%s=|J�t�T�C�w%Ùގ���z���:��e����銐k������`���ʆ��fD�+9��ʶ&I���v<�y�,��m�B,�C3�`eo��s���'_���r�>E�Q*� �����?��r��i�:�̊�m:�ￓcu�����M�?��t.'�!t�s �ֻv���Rn�̃���[WM1�$��GU��n�޾ىok5����h�������0`�(�Oυ��`���k�%���!�`ܧ�j�l��F���#�z�gE��6����|��Z_��h���%R[.�	z���)!����"�[&�Д���A\��� C�`_�F�2`�����^G�����O*Myo�������^΅a�>���b�u������;����i��'d��f�}��wh
���癭N��o�Z=wQ���F�2""�f2���EY-U���s}�fs��ո��-Z�����`�����9!5��pYz(J��0��6^g��[��,)�-��d�1WE⾱��N��S�����ӿ�0
fU�j��+�� +�4���z�l{��M��y�>(�Dr��c�=�42=}G�� M��E�>}�he��Ve�JƛjI�]87v�O�������g�����Yx�����#��?W�l={��e�D�)XgT��#�d���FW#��J
)I��􂊘'$D�����H4ltTH�e��^�X�%�����n3�M��w����� 3�j���WP��Sv�_�	\����uBP��1U��U��A��D!��n}?\8 ��^�?����Zw|"I�+�֎�"J�/�i���9If��/��p��b+���(����ː�%��#{u���Y�GX��$qh=����Q'���0' �����Zo�)tܠ�	�ɖ�*�g��w&'dԣ�m��wi)}�&p���1�Uf���2��[���O���9��ͥ"���WS9b6ڻ����z:�v�g������X3�i����p�V�}[6���{�;��������z���1�U�>ch}ܠ�.8��+I��:䴑�d	���%�p↽�yI�\9��.��X�!ws��X;f�;�Y����|0�-i�w*��P|$
2FI�����lA�PH�*��� �7�r^��#U��P�NsrP�ąt9;ɂd��h�����,�Hg>���׫�m�{P��m�a߅������Y�q �xzѷ?�F�EM�>JD�~_`�Sh��c��B���;�׽Q��S��
2N��x��(�2;�.�M�K�L;�_.�#w;t�z����lڇ�1^�mc�{k��&�$�<���#G�n �l���e�|s�>��ۨt�w?=9ޜ�Tb��l{}�6�_	��U�k�h_�B�CJL���Q0�i5_�d�wH"�J�Y�k�&W7:��:��g�og��YШ�ڮ(??�nt2�����{��T�$�dP��֚������Td1�{ �L�0�GE�\f[�g��Rn,VH��:�!LΈ�D�]_ULL,nb�����j	]���Md�Dg����;4�O�q �{�)¦��;;;��]yY�B��6�qU�G�3�2)6�ç�}	�FcS)Y_^Rc��뗽�%GR��6i�մ�Pye�"�3�.�E����P+V"����^K���������ɱ�
 �ex����;�vO��.�Gzt�l-��)�����X|�"�-V�V���|V̩���������R���%�j�����)�'�񂕭��@��=a��Z��+�&����?������	H6��,[�[��d]���h�OLL�ߺu��y���9�_�#߅������*�<v-7��^��jC�3��(n�e�k�w6�N5����͒:��8�XN�φƈ~�wj_7��LȮ�Έ�]�>ݲ�v��K�w<��`�(MP������\TG�2U��5f����QTB���%��B��H�m�t$^p�������_�06���R�Y�����gf����J/<�qS��Q��rM	��/F���4�B_���+���xu��p�]@I��՗��ȯ�o@�RA7a�C?��#p�.����kc���>��>Z)�Ge+�2|ɡ������:tC�')ULg�T�@{G`����{Q�<@ ���6�T�� ��R��v{��oB�-�3>S���s$�,Um��4�:��+b�C�B�nwu�/Ե
C�% ���j��|��g�G���L�}V�
�e�l&;; �-���
ލZ�������D����zIƝ�|�d� �||�#Ŵ3��qY���������-Z�M9�� eF+-v��[��Q�G��(�Ł��z�����|���M�>��|or��W�f�،xW����զ���D��0�S�A����lS o��}�V��mٛ��b0��8Dk��C JH�<A#AQ�S��U� ����8��>u!n�ۢ���7�4����|W�i�t�\;&�w[�!���*v�wp�x��޼{��Y�/�g�:N�s
��=��$&���f���IK�������ӳFG)�Q*�c�%�ˇ. BM�?m�����*�GG$�Tw��o��q�0����M��ˢe�ư����3��������ΖTj��6+3R5�RϔfP���74ƶ���0j�W�f):���R��S���vJY��3�@��nQqޘ �ݛ��tYv�77�y�����[|�e�IZ��U� _X�e\i\���$�\gyi��I�r\��ӿk'�%vyj���S����C�W��֑��R9�a��|��K�΋�Y�RV������c\]�n�@�I1���D�e${l>+�'�d�4�_����B�-�;飤t�D��ؓA+���o"�̠��V��ר�m���nj�]�nl�k,�P �7z	��H��Ho\=B����h��Gbw��l!���V�~�s2��6���ۻ��D�Yo�p0y���+[l�T�
|N1��'ίѦЋ*;��xD�u�-�'Ľ��Yht�]U�t ��@��������o�8z�!�IF��:i<$�Sq�4�9��ʱd��a[�
�x�#<_�%�F=�zp��̭��:��@�^��%�~
�m�[�ō����N���Q�L2r�MD��yN�Vd���|@�,��?�ip�W��%�o3>��C��L�*~�D�Tc��9��!��+vd%<��O��;.b�$�D���3�<q�����Sf͍^�������W���k��"D�~��VoKO=��z���B��#�='�H`�q/
�Q��Q���Q�A�`��v3?j}���h���Y,�b�KW��������gP�$YL7�������ۣ��,
�i���w�C��\^���,��qf(�T�xP����]{F]����*��1��XQT�?i��ʭƲA B�-n
;d.O>�*�	�@�Տgp�+Y�銁\K\m6>�Q���g���ۧw�^���4̄]{3����:@+1���r��i��>Bt�����f�I@ʌt�Y��a:�Z$˳��c�]D<��g���i
�6����Z��W�F1C�R�6*ߖN�3�.�P-�?!W�z�`�Ü�ʽ�Fu^`$����&�ʃti_��6����`ؕ�Z9�7+ *3��X�����HU<����X� ZQ	U�ӳl<.�{��$-��������ob�L��S<���VΒ^�YTg�N��;�ZO�c�ם%�>�i�*aľP�)��5�4�&n�<�W'�!p��A�)8�gmm]b�8/4(��o����b:�td�W	[~�Y$��������9(�TJ~��I�iPYub�u�6Ӡ�(Í�Wt�@r3�6:�kw��.A���'0���sB���9��m	�Xn�t����R��Ԉ�(�uzsf�,o�:�u��Z\�\���Zْ����!��V�z��©�.d���S,0f}ԥ7���^����~���i��5�p�#c�Z����(#U�AF��t���K�`�h
���8�]�c�k�߄�):�4����q�F�`����i27#�����Ɋ�PضG��P.DbtHH���2>�UK1½LĎka�~�t�UV�]��3O�q�sy8E�߽=�+`9�����!��͟L�Y�ڧ������q!VrZ���M1r��oM���i`�+J�]%�5���}�� �ԃpf``�FH␄6p�]-���23���Hw�~5�������v�V��$�x��A|�L�-�l�Ь�wn:�b�w�e.(X����}b��}���X|�wW,7���w��[�}�{���5�*�g\(g�E��>!B/��o����/���Xڮ��]�DPzw_8@��>Kx�&�Ѧ"K6���/��@�K���ó��X��)��獣:�#,�1,��j����;��)(���MJ�����uP�7�[T4@��Ï���^~ڦ�S��Å�����b��(Mb���~8z��s[�ʬ�{���S�4xzt�ƫ�=թw���Q�w�����콷;a��5a]q�`�]�VlOG�2���%145���{4u���S�b�Q�Du�jar\o�H�8��C58t����"ˬH$o%�{4sB�b�J�*��cH�u|�y�F�Vc��e/� ���V+fb��ݕ aW;[Gu��h�z��G���y	��	��&i�ӊ fr ���ߌ8[x����[X�	NîsN`��W"Ia-�tQﯶ=�\�M1ٺ�[ӳ����ݬ���T�A>��*�mur"����oPL�U!�cn	�s��~ybC�����Bǎ5/�o����v-�����L=c����e�`eȇ��[�z�l��ě����u�fn�~٧a�%�f�J~c�_�q��0���>��SVt���P�2�Tq�Lq�P��?��^�#K��=ZsI*�v
R/k�~���qB�;N��������1r��.�͚��)^&@���P�x:�p9�@��R���}ԫ�D�ymIF�BL��������RǕ�d� �J�5֥��̹{����I��{�v%�\��eo�j��r���a*�`�\V�
t!_6����j���ԯ������O���l��X�Gh�R�1���R'��
6��[�n�p��<#F�N6W�xe��7����C��NĄ�I[���X�XB�몰�5ٞh4����R�=��V�����$�ɗ*�����K']�=��=���My�*���/ONV9f1I�����c�o�K�*�>}���/�|0��X�K��
6������5��#U���rs+�8�E��B,��֏��J�9���"(ب�۫֫�L/&�w~f	���|��U��kK';E
#��t����e@�skDv��'�F�}����o��/&�B>��5�A��1�oҳ��p�/��{�����?��+<�'A[5:����D�<���]b;㥽��	yV������{E���JQ�e	y��w8|}oW�2@�c
��[��x8�k�N\*���!Ʊ�7iY�����_ã/���?��qh�栩}��n�����.�{�I"t����?���ɉ����4�?�B�b:��������c�y�R%����2�M�oS����/�\�p9�p�I�b�}]�I�3�!���8�nG���Q���޻k���LU%˾��߭6*����}+4�'�zX	ò�b�[���k�QTa���8��i�#����7Eu,o��� +mP���]���,��Y�m����c��w�:�����#~r#<j,!�j�t�������*��8���Y6Ҽ��$OeP�@��<<r�M����c�AwM{�/G���#3U�ķKy��<^�p���Ehd<�3"�죴�u�E*V�������� ���}b�;���M��Q2�s�ɋrpD��h]�s�8��wb&f��_u�JM�W���3��5�P4�tQ���J��=���kϱ�٭g�nE.�-ּ�P_mʻ�I�"�M�e��Bn��(��w�	��Υ��c�����$�7*��F>�\����Ɖ	�)�x9�͌&m�R3�] �����H��,Y�r���w{8������zo��3\;�)2go���:.�j��D`��2�{a�w�r��Lets�r���rw���V@�z��y�y#�C��5�bػ\����x�����2���2M�E	���ҙ�hYݱ���eާ^c�LBJW�f��t�׷��M�m3���|4/�qg꜏���v0��n����*Z�1^�B�E��Ñ�MW��(��ʿ?�Vv����F�F�(V�V�`_U*�����;��1J��^*��+y���=��kq�-ԯ1툸L~�W¹8V���)��0$`3Y�Vl�>m��ag#r!X����~i�g�Wٽ�����/��HI��9����7��Ŷ)�~U�O�61RL�}X��u�I%��2kٴ��R���\:��b��_�Ӯ˓��T�9��O"S��'����Zy����?ڿ�˭���u�*'�9)$�%Y��J
��f�D�������K��"�H�e=@���z��×�$ױ���E�_�3]\�n�ccl[=jQr���Y�ȰM�]��R�,�.��ׄ������G
![�%+N^��/D_��A�&W`P��W�&<3/��L�<~协�F�K� s� d˾*��Lu����<�~����K�Ry=��~+������ྀ���Ƀ�k�8�W��>>R@�O��rY	[�/t�3��#�!�9=Rnyh�X�� :^��bf'Y�M`%�mkWq&�ѹ�===Ɨ�Ih�ã��G��������c��o(wAo�l���3';U�������Nʓ`�(r�i�4'��K
w�,�IA���(4h{�� �!��>*�z"j�.��.�0Y�覇[eƍ�.�ׯ_�v�E�.�m1+���p0���,�Xn�e����98Ȼ�Y�	����vHe@&��6���]|��v��y(�����DPB)�"?�a�h���,���?�:�A!�7�s��5�%�?W���K��W�O�0�V�x{�s�gϞ��A���4��}��]=����K2�nCVV�RY����H, �����h)��.�i��L�G�k�[���?@@�ܓ;l�z�R�����2r'/.Y�[O�����aQJ^��x��z>E�
y��z�">�:�q�5}Û��4[�\۫r�[�?�<ݲX��s7���H;7�gg�S��k�O���g��4y��W$�i?~�~�G�ҫ��$��u�D��[�%��<�<�<�I����Tv���!�������#@~�DE����Гp�s坹���<�V	{�:h&���:� �̜ѓy0_�s�lO���Ԯ7����	^��A�6���$��[�+�9P�!��k�5ZN�%�y�I��{Ue���2�� zE�ܕ�������	ѽ"��%���9���O{y,���k~TT��t|S���ɕ�Ҭ�����	R*8���Z�����	�3������^̉H��s;,ē-i���V�{��@�b\��Uz��وu���.�t)3�T�-@B(��\������4���M>'� F�/_���Z�@��J���-�LU���j�I�y�� 'i��0�Y!Ǚ�����v���[��!������|?e|�@U�B���7���ڂ:���VS�UY�~+��)�1�o����d1]���9ܳ窇�F?�q��2]�["~��犔x
Y�N?�� �����}B-�Ғ0�����'zc?��H?[9]br���,�"�P>�7{��_J�C �aH%�k^�}�׌��T~�۟�Id�f���)I�3�//x3��gExX9��^��s��ś�
T�U�/Ɨ ��~ދ����M�c��w�mg���5���c��x�	��l�%M�s�#��w츂��rK�{��n�H9����|�GRL50��;ܖ��Ol��]��Cڼ}�ɷ�p�������gv^dv5ΫU ������7E�r�G�������]�\���E��0-��PE�k�o3n�p>�$m���|�P�#�m_ͤ�m�< o7���O��(7��W��u;1��'G�Ie��Z��更`��)��|����%��W�e2�O6q��A^�p�.�6(�W��ܙ��|����[��Õ������Oo5Z��?�K-v�ظ�2�t�a�Bܗh�t�]���}�"�/y�vg���� �v�/*����k��3��zSh�L��*t����y��]O���Ϭ��q-��$��2�(��:�T��ɋ�`�we��"���0D��9ي�1]}	}bG�n��A*B�L��>�ΰ���,�׎��$5B�+���U均�1�>׎^�:�AO��L~P�L�C����/A_V��ƪ�W��0*���U2����fed@�~������はM�3���2`$�`�������Ŧ#t5�fc�~�W���ϧ������L��)V�<�%BS&v!�����Z�z��yf��������=%ѝ�t)��!��b��;���X9�,���z����R0R�5�U�k�'���|'�	��C���a����h����w�n^��eM��<9>���}�����M���aA ���H��|�s�3u���s.Nh���u�)x��D��yO�]&� ��

*|��	�AŮ��\<�؋>B_��ZLL�V/�,����*������|����1�5Q�#��IF���S����P=��o� Eb��+�+�|�,���n����ԍdD����c�ԁ���;�]����y*c9*S�X�]�*S�%��d(�2ce��R^NfU4QYZZb6[�Ӏ����U:n����go�.�=��6x��r@�=_��g��CO_�*�Q�g`����B�X۟H�[ڜ	kfd�@ީrǂ�w��r��8$[��K.`	c����Du���_HE�^<�i�fӉ�\Q�0��Dc[��Z�`����:L���W\���Z���Iz�CɼqϏC+��M�>ۂ����؁�Ne�j"Ǻf�#񚆞�Å���nk)ޢ���Px����hd���Y��~�'��r�^����<��l�V�5�U.EPB Mm��%�o�~C��A:#B�
�P�������0�_��ua�@� �d���
���QRd���%�3��'n�s�8]K�T�0���W�OX6�I���6ѹ=������hټh�I��KS�9|�<#�3hN�:Z嘃��|� ذ(R꼪�]���o����bF ꖗ[��.��+x�Ho��|�U-�V�+��.�d ���F��� �	�#A[SR�g����@U�!���\�H1Iv�ho-��!�i@@L�k�U�<��8�J��n/��[�c�ECx���  �����WJ��������X�cz��O8�#��-6U�@V��뫶����|P���y#��t�>�����X�3ˬ�uy\5�\��J)QH��lwo��,�P~,��χ�|���&��(qIO����uN����m�Ήr�v�r�>}Ϯ���!0D�9��DhFƛ�������0�!�V�����/�{{��.�{M`aaFc[���MVe� �4�=�V'l�]\{����w ���E��t�楿/:j�d0���*��Ց�8?]�� �c]�&��ҺB�n1L����y�[ރ�]�Lx���tжŰ�-��pee%�`�!�I0�����,��k��1@���;ڿqM�K�����C���8�4I?��L���� �� �_�w��n� ��9n*�oN:*׼���k�)�չo��>���1I���d��������ggk"@^�	̯�7S5]1��.�k�]�������gN�O���gĄ;���^���
 G�bkGE�f�
�?D�"�&@ُ:ۉ��më,t�c̀&������� q��T%����X�ݭK��n���LT�O��jyFCL:�|�]7��|UC�q���St�b ��ul��j���z������y6�:
�x����E�?��2k���
'l}� �Y�26Ӊ�|���?���Sv�t<T1�HU5h�-�ߋ�a<��[��T[������y7��S���y�H����4)׸����8��j��,�gI�%N�2��1F6����9��Kt��t�.��Ժ:�(Ŏ
� 9��[!_�7Lw!W�T�$���^|����߃���Ͷ;3��J�u�$ 5����Ą�>��ޔ����@���� =�ǭ���RU� ��QT�|���	�T<T�JO��m/C-��d���f�'���z���Y�ߢ�C-��d	�G���#��˔�hDDL[�Ug����,��~Wױ����?]�2#K���2��Ʃ]Ȫ�f�ɝ��)��&�M����,U�e�#���]5G>RH�V��P����|����*l��=��U��� )/�W�q��]�0�oh9���� R8���^���b���y�)���/h��r\Q�f�pG�'�,2ml��=*Ma���m������
A��d,,�r;���#��~6������(�˰�)��]&������d�|�G�ʽ�Y ���{3Egz3-l˯H�v��+�K-�w���b���(-�u�A!*�D���m�{`�1�u���1wP���W���r��'~V�P3�F����<7�O���,���T�H챫܏f��{&�E58������Cp�ſ�-(�D��w�G��S<�E�j�5����I	ob(B�����RV삢e�o���B`RB�`�^]%V�H	 _>�m�����͛�v�kv��u���h��j8��\�YH���Y���-�������CU�>�TVT��j����l�w��*?H��>��L=����+�"p�����>����p���Ϟb�^ �%�>{���0�۫��\���۴�%�2�#@�0��C%�j�������J�M^p�me'�����/����'��F��bzI$�6xZ��������	p�����q�M�+Z=l�ʄ�c�<X���.�$U��r��+�����@�L�����
@�F��Dr�^RwS�[])8rw�NT+{4hQ웛]<���n� ��z�}�2�ϳ!�l� ��$���K
	�9p�%���8\��(g�7b*{�e?���tL���u�*䴆�d%p9�����;���\�o{�vhӔhH�
�˴�ֳ3�(�F.9�z��M.Sf��s~O��Z��?�it��J=[�6�]�~-|�f��v�>��o��%nb:J�{{���/��\���%n�Z����w���?T��9�;#��z�9�ve>R�y@l���g�˿��<ff���t;�{RL'Q��$��E$t��?#������ȹ�rP��RƂ���SȊ�>�+��+R;5J A#4��1㔏�5w�~+�]�=Z�em�8$��z1��X4]���b�8Q��d#(B�t���3�S�����v����s��4<vì�BЏ�N�.�jҟ����6��Q��ܯ�4Ⱥtt��;�.�\�ڭЕ����J��=xHb� �����c� ��J��@����b�w�ݨ�u��7<�+��dM}Q-c�~8�	�r�aTT�z����Ԛ�����̃�)	��~��l�L	-���S��� �ާ�w�S���������M�<X ��Ja1RIE��-�k(�5XZز�|�O�K�����dR��] )� R�ja�f�)��Eqٛ�N��c]qm�n~)�P���(}�ݸ�D����÷�+�z>�P���_X�KS=�M�6�fN�A1�j�l�@+�)�4X�kkk��v̒D�L��������3��:u@���nzk��צ�B�x4 �ǘu| c�)�T< �%%tC�8󉎰#����4��5�)�G�s���9��&b$C�BF=vC� ���2�_���U#��[�Y�JG��@e�������yOpƣ{o}a��a�u��"�:��L@ ����U�ޑS9��Gυ$���4�����3�,��X��1����~�Zu:@�6��#�

z6v����a�$;V����AL�ݲ��-{���B�˿9���)�u�K��A%`�eBi�p�H��� 곲�z�c��
"1ו M\�����<*J�\i���$��AǨ�x������dПw���V@�͡��!`:8>Ξ�Q𛮙v�¢�񵍍F��'�:�?�#@�蝴���đĉΑϹ��Rl�=ޫ�)�${�<��<�����b��? ��If|V5��?V54,b���
�����l��e�ʌ[u�K���I7y�s�Z�b����i��7-��PB���C|�lD^���|̍����OFhD�h1�@�H*�%U��/.�Ł�4b
���������V�@ʬz|�	���N��{C�@��Z��'4P�7��pH�
R�� �>=�-�d�n�Z}?v�/��,dYo�f�2��&�)�y)/2���0:�2�ӿ~�2���}C_V/��?�.��R��K�����Y�3��{aw���9�j,_ߣ��Bw<��\>��W��E �`�,Xﻓ�v���.�N�[�1�����������X���)t�sX�0h=�#�L���������OD?�hFn) �Zʭ���&5u?/{3/�p�	083�aT�#&vqPR� )q_?��m�`�iH�<����*ya�jߺ��8`)���H�=ʀ�7��� ���&A;��,4[? q�R�;�7���o~S�.U��`��Q������o��
�K��t
�
�\i�ːJ �qe)a=���5�����&�K��j g�2S���/~(wk�p��@�v��
��%�!����a�n^ �T@�%Sd�^�f���s^	C%�?Wa<�|�j�ov�Aӑ��8c\�Z�9v�-�X�̺�PƆ�R�0%��8U��{w��П�F�b����0�����p#IhE����/JHI��b�+l��� ��
�t��T����8��[P��LU/b�KR�C1i�X�&��}Ƌ��)��w�a�a돤6�F��Ԥ#���xu�x�v�k�r3y�{������$+�X�1�c�jڇ5=�6�r��t}	4�mԶ���@B�B�P�y.S"�p����<dh"N$3!�1T8f*���9�c���?�8�����[�]�w����}�{_�������K�2CU�����b�d���-L�0�^]��Ax��庩S�'�!J ��J	$�Z'��'b�5p��k:@�ɣ��B�+~]�Y�4�J�x��c �!�u�T/���c�������A������C&3�n0������rO���x�t~��G�%[�.,�#j�]8�t|��٤r�?��ʉc�>��:ـ��w,��<A@X#���>��_�r`���w�	���Ue�F�څP�i��W�U��?��'��N%�D\!A���|��5)2���`���*wSA>���~�4�	bS��N���C�A����T�+_N,mSgh'��q��FM䩼���a\~W�a�_��ۉ�������J����"��;�9g�vaq<O�4uͩl��bl�mhb"tCF��{�Lj�c-,,h��3XsTw���"C���_��r�Rg�����Գ��?��V�Fi@z{��}y��,��f��ͩ�r5ޘ'ŦXRA���%�sl۵K u�vV���I�"�¥q���O��V�噀d��:ϔ�/C8U�f�ѧܪ7�Sf=�11������j3�N���k��8��C�6
i�R��BA�r�^�:O��RQ�!���q�i ���B�k��!��@8x�a?m@ �	���K*@AH%�U͖"\�FV�ѨI�̄��B�`��w���D����W�	�=g|J��U�;����{�_C)���W�`7D�|��Kp��{tQ�!�9$34�5{�mG���5�os�RO��.�#��Z�3��D������	t�aӧyy$ʄ
p/����b^l��L
{�/t�P���S�}4�����מ8�ckX���)�Z�Br~>�S�K�kC��4ueF��j��+-�8�O��;ߺ��@:�z���ݻ����V[N�i�I��#]����LϨ�CsQ���f�*��;���f~��N逺&�V^H��D�Kp`�>d_���_�7�Ib�b���-x
� �h+�E�9H�.�iE݁@ɻ��Gǻ	q�E���(Βêt�/,��O��G��Mg\�>��}'O=��UR���3f�S|322���Z�S+^0��(��ڴ�oP��$:�M�ģ�	V*e �)�@��,��`��|djsF&~�#��\b)6z�ށ����꾩�v�A�4�<mp@�o��(5�vAE=� ���r��Ⱦ��3㝂(;����w��hI ��u�C��rL��,v��� o�
�=A8�>�j����M���	R��ڬ�f�*^�+V)C���)X�rH�q�	�����| J5�Ρ�W�*fg��P��R����Q^����Ry��qq���r�!��lV���O+;�d�$�"��5�Z�o��~$�hTѓ�Mf.\dW}�@p$f��Zd�W�g3߸޺pjh��b2tZ���;d��+���� GpvnAv�'�iC:�z�<vL�Y���;��iL�3����wA�ֺ�/Vw��2�W-�Jҹ.I�����`n�}�Էu<�	��2�S��3�/��S�jQ�����ʭ���_�(�50�27#H���4�ԉCj]*xd��=�N�qZ^S�(� �6�� ���%#i�q�JS\A#�Nr�BpW)�4�K�֥W�/4����4Vݤ�޶��?�Cc�W�;�\b���ٯ9��ߡ�ڋ�%-�����/�P@�3��6���™ѵ�i7v�IާCv1|se��r��x�q�ImE[������;�1Aq��I"j�u,Q���U�@�T��3?qi�5��Zj���y��ẓ�-���٨ �U������v�������ƥ7k�2f�ب��MG�S�~�E��'�}O�Hu��pJ��%g� } 2��w�1`�X���������¯yrW�+#%^䨦p![��CۈWc:c�빶�ըٴ�	t~_�шw��A���u*Rh����>�)�Z��[���E9)Γ�>={�������G�O�n/\_1�^�Y�!��KA���������N��gk����iyb��o�(�?@m"���O1ہ������Z�lǆ�7�}X�GCL��<��Ŝ*�*�DKvp�m���zy�X�xj���z�"��z��66619iF8zK{�a���V���G�P��=�2�ۻ3D�	t�`�A�;��S:k���~<�6+��sD Q�WB!���])ר�J�$�ɒ8n�zh���a(2���P�:�����;���(�Ly������R��G�5�G˖U���)[(k�`�c�.���?���ϯ��퇲/�\�hK��/���6�?��2Z�U ��������g���O�5)�����C�^u�V�x5���I91t�>y�$G�g�M�o�}# ��P��n�!�S���as�O-i���l��S�C
4#����J-��o���!���>�s�[	���"�s�o4��K=sV��6v�?{z|���]��w�;'����xļƬ���[��83	��)�s�����N'XS��*ʊi����n=�cO�d��-{�#3��6R�6��.}�YB�^�w��&b���0�Y�B��Zf��<���:7$G�|��+�k���Q�eYԭ]���t��?ud<
˒��XM�	W�{�8�����讆ٿg�0n��5�q0�N��z��X�w�=�r5�7I?�+�������G�6�1f�;(��A	���AY�@"���_�7iJ�|PypY�Ro_���G��2�8}Ӯ����`��8����H�vܔ�
��k+M3����� �m��L�E`L��A����7��P��9����/u���-��]���{)���p�SF~ڬ�aR�Aμ"�^�T/�^��q�qt?��ha�9Gݣya�v���q�р�C���鳡꛳��,g:%�^�Rלh�����1�4	����|�(e�p��7v���i!��S�y����5�}��;�l��[����>Fh�Yխ���u���fN�	�U0'����>{+-&-���T޼X�n�蔴��I��<
�����8�O��/�HD8��Q�Zk��2c��/��������0?��%� ��wM�fB|��*մK�g@���{�	�:�RJ;1��?)	��u����<Y��#k���s��;�@��!Gai������9`�V�������L��ʣ�#`����[P��O֙9-�Ͽګ\"��T�����N u����U��֝W�.���N�L�J��1R��y"\ �9���*�W���9���cf߮*�Z����,pڞjF��������τ���2��k�!��i�����߸ ��W&��c|�@�U͟RQ~��T��1��l�Yq�+Ρ����҅�Ҟ{6}���x�������t���|E؄�+w�L��DQ^�?Z?F�)zX��m�5揰hp�6��:��|e�*�b�j��[cmQ��R�I)����y���Bâ���~�"#no�=^�
4c?"���;���3��C����7��0u
v�}�Dg���@�r��p��vw̤%��6c|t�Y�R��2J�Ϗ���S=99�ő9�"���}��吹˥?�\� �9/V���KH@h����\��5j�܏М@Z�@?G�R��+���Ԣ?o4�ff)e`�Cv o�F.�h�*�T�����J��t|���@BL�~�/P�f�����hVZ��ly�V�_�;O(��̋j7�dk��`���N0J���;~'n��ḨG���3����)��O+���=ڪ��ѧ��G��Xo+/b�	�.�m�OD��Rr�;E��؆O`o>q�Έ`�Nr����%�����qo�E���j��Ɛ>m�B���C��3.,J\ s�7���x�N���E��w�V���T$Jt�p�ڀ/��{*�������^F��<�+hx�$�9��E3���a�d<�ʆ����e�B[o��D�Ѯ�����ֲ���ן6/jTF���2��Og��~xU�_58��e݂�ލ����F��ٖ��y�7,^#�����Nk��(֞"����026���[]���D0~�(�<�S���A�z���@�{(�uP]���@)���JN}�L[�!̚

O�.?�S2p2�$KǄ7*	���K��$��,)�Y�W�;R
@f>5�n{��}��+מ�
�#��T�椸lǉ�����1w^{ 3;4�
t�9����$z��?��Uԭ��՚�����L[�v�_�VV|6T�G�&�8�K���{�CԓE���c+ ���\}�������Q�8���*z���T�W���:_]����~&$C�o�v�Ģ��d�4fd�T���o�dpl�3�K�Ɉ�~����N�_  o)�������K�	�g��KJEQ���<˫ �����M�=�+���hk)<�'���g�׶�$�gk��,S�s[��!������w3[�&TI�h�*��&�y<=#$eY�F?�L]�/�':q
��b���ۿ�!ǊXo�s��k7]�0(�?�q;3�Ϊ9��.��=f\Ą���V��,d�jm
 ���1f�I�����;52=Fwg� C�/�Cc3���C�H�UB�#@л�ol����֌k�\�9�Ty/����ܭ�,��B
͑�z(|Y�R��\uBc��GE
�<F�(�&��*�eۯф�j9e$��$�sGz�K�/����	Ks����՚_�Nb��	bN��%'���Ӣ.O�߹��!��kʖ�=��I������~	6Z1���ABq�Y7��������5"DBO�ӳ"�����S�ІOKa�31c�c��$ �Hٗ>BX�?�v��+�?��Z��EF5�"E �z�m3>��Ψo1�?�u!��m�[�lqv�l�]�ym��"�4�`�E&���X=�0w��� �X1����
YGaS7������?[�r@N��Tf��(�oI�ǫ̫�o�f32�2�_�xj�����6ѓ#����⫴0+
>!���"D�T������f:A�G��ޖX����ݧG���\�����S�)�b��9̙���o[�E���Ƙ%3 7��1d�)))1L�66��Pby���h�Q�ؘ���c�tAT����C��&�:>WT+[t�˫�G�^�@����.?��0;��������?ߚ����P� �1K�9@�Ҝ���o-�&�p&H;R�&N���UuҨ��1�]�� &UrPt���Y[ �w��4�����2���2�/(�������+���c�������F���^��a�r�C,��
����13s�T��TZ[�����#��M�D���Q�����vv������g�^��?K���du3�����#�[4Dr���%w��,bG�����I�~�=�ؗ�G
H�9��C��|���r+4J-{y��.�B7L�����6u�Zz�ˈk���l|o~<~-��t�����?�3L�5���D�n�uZ������N��k��u;�z��V`߳��R:g��4 ��1!��j����{�N��6�$U�����Cv�m �������� ]�/�Bad)��V���d�w���*r��*�M���1�v�m���% ���Uk����`��&T�%z��M��G�I�fF��&�x^X8�y���Zr��x\>hr�*�$�{TW�R5��3�f��f!"E��$�Ǳ�#c��(�2�SBC�$<�������`�%�L~yjw�$:7J���5Vi4a������m�uVG�O�z�̨�'�Rs@̂D�.<�H�XSzy�����f���2o�a�Σ�+���J�6ݖY*�%_�D�D�4�2���O��%�e�lq/����r�����S�k�M7{?�`+��.���n�3�w��oaDX��Ǵr�V���ܦH%y�x5x�P;���`��766Z-��Wl��s�?�Mϸ ��D��q����C�>j���/60���in,z�߽��3U�d�2�<}�f&C�)�����5=VBfH��k>F> 80�j��	}���@T�#�u��J�Y�3!�@�!,�Յ��c�>'�{�Mh|eQUzW�$o�5)QM0A��O����� �=�m�_��v����u��p� Z0�����h�~���6:��_�(Q8��n�Ɔ ��)��Dɺ�]9��ok���FS��mӓ~�Wrd�c�Z�0�g��s���g�v�e#r�Y�a�v�ٍ��L$ҐE)���}H2�];����\���޿d��hn�E�Ѩ�UW���Fj`��c��$Lz��ww�*b����2�Wͱ3$9�.���+���Ϯ�[�QK�iyzbZ�/�:.
_S�^��h9��P>��X�3�}r�<��8}��G\	&��1K$K���s�y�?���'�l���9gAV�:)�-m���کKScR>g��#��)�,�<߭O���pJwB~Iq�rAQy�t{���;
=���<�㼯Z₸��D�ZFUzdǭ˃�Y�<����j�w�WȲγd!\�g%��v��SMd|��Γ׬G���x���,�%������Qg��IO��N!:��H�-�peͰ��	#$�R�K����b����[A���j
��_.���Į��+Czb�R1`|^ '��,yh�h]((,{A!��49X@��C|������y|�;u�oE�~-��8fǱ�OT���^���������"�q\^��x/����{�lc�Vg&���5�p����5b��y��Z�W��Jg[���3kUSo�L�pHK�'{���O��T5�G����!��N�E�9^�q�R��TM��kB����C�W�	cX���g����r�Z���
�p�۳�s�y��(������$n��gJ��>]�G�B&|�QVNY�P�,��R�ڛiF·�痆��s:��]Nvx�T�ѫ6Ad���ס}����ף�s���}�fr>w�/��u��� �5R�l�3�-D�L����'WkiT�+;bBG�=�3����p��=/�#��D(4�9�5�_�;sV��o�����O�a!wO9���޽��[+�f���M�`���[p�X=�Te����Gll�afdD��"�ѱ�7N��E_S�q"�������v@r�oU�V��Y�o˧C���B$^?W�"��^��.�m�=9���j�.�W5őJ$���:΍�no�]������lF�OFi?���a-�-3�$ ��Gaj2��CB|mI3TH���_ɇ�^"��H��{�n���G�����O��A���m�Q�����P��M�odYHp��g�\�Z��D!��,�2�I����H!���?Q�Q�*-�m�w`�1��5�Ͽ{�տ����E�x�v��I���H�(4�NfS��9+d�nIi<K�.���f>�ʏ��G�1�#��A��Q���O�����8j�y诵}!'}��)�g���X#D��H$wN�����T�!�kܤ��&G5�er��&+�� ��>Z#� `r8�S;�.W���o���Ӝ)&k2� ���z�&XCT�_�B�J�H]�m7k���Exݼ�"�������\3�V�Q.��Xٲ}���I:w��Ї.3_U����$�|�w!���
pʿ���O�[}5ꅢ27k|�z�ȗA�ƪ��q��b�|�L9Iq.碆�}rr��4����}��$l���Qy�(*K,%к*�a�ڨv� �E�s��H��PW�SP4%k�5�Du�<��Yw�xqRcc/H냙��F�7]�񪫫�Ix:/���kh�S���8>Q|���>�z���+�d⽾�V�ȟFvy+Yon��@���g2_�j��M��g9��[�[.}�u���'"&�O�V����n2x��1r��e����u7!r<��3�����d��~/7���hV}�`�$�����!�Nr��*��#�����iU'
|X�M".�B%���ǆ?�29�+;J�[�aN� �G����dY�D<S����{�yr�L��'� �ld�T�Ϙ�o���T|�ݣ*þ����9K���@GI���3*H�5�Xf1�F�x�mb�v|�B�@@5�>�Z�D]�����r�3���q24�&��\{$p���[�$��IU�#��̷��m��(q�A�r�L��ީ��Nb0e�R���Jm�RH	+98a#{Vj��v s �ǈ��\lHTNn�|]=�2y{��0��쒁�E{5|щG��������*8��b�bڞ"W|f?�P�/"E�mX�Y�S�L���T��J�J�$�-���6�l�;��q�� h*�B���9C����z�U�fԸ2s
/�[
�C��Z�'ʤ9�{�u�s|��f\�ڴ�µ��	5U����V*�	���]c2 ��EB�Y��@{����X/�Y}�9�.؃��1|�8Y��f�f���h��ѷ:�4R�����9զ�h��B�؈0��K��L�s]Fو<���$��v���S,����X���uaa��Ԓ�v��1�F�[A
�L��N��2[�a���͗f:_n�([�1��p 9K|���܊
�p��<����:���݃D#�dL��#.�@�w�������4�zY'�@Q3��- !��\|�A��Y��_����Q�4᫷�	c~3gǍ��M���h��@�ن�� ?����fF�c?����邡k|
�ʄ���S�y�ACuu��K��3�E��P����e���������$�2I�\T�_9φ7���I�2u�TV0��V&�rLi��&��Bz)L�b?l���'k��'dyܱ��)�9hیJN�&�>o��
|��m�a����B�\k���i��j:�>�ʀ(���^�R�bS���,���a�|hh"p@����?����sO�e(�A:E��:?�V�\�!)�-�pE�l�!����r��h�
�4s��m<􌿖k�5������,�<�9XT�X#0�b�����f�&����rvalk��
:�O�:�q�4�3�! ߌc�믵����|Gǿ W5��!�%���S��XJB����q
JA��q���j���B Jo�O���V�5��a���1����K�Pb������Fµm�&����\N>_PoU�������G��C|{��"�^�D��۳����P��P�xU.��F_�#O>�.���q����"cO�������� �u����}�RŜ,Bʖ׷_�D��O�y~!��S{��T'�w�mŶ���LT=Q���Z�z�:�sts����4��5 F�W��aj|�Ȟ��'�O��F$��E�sf8Y:��`n妷,��nL!8����g�?'��¹�z��,u�u���g�n�n����7T��Ӆ��x���<�xU~6t��^��g�^)���Mr�CIpb�k�Q)+n��|�ʳ8�Y���H3m'�"�,��~��D���/�s*�S}d���A�����Z��|�����s��������3�B_@��5+wl�F�����Z9[K���q�� )��M�!����l!z�|BB�m�(w|q����n�#	5:4p\=C+jp���w�ښ�7�_�sx���w�#ђN���]Y?%�4������Lsiz�m���W������u#\��A:)|� %m��7�|��ZEq���뤷>�#�5���pB\69J��KHDD������\��5n�V�~�7��lUq�c���S};D��{�&�����������WAb��gT^ńz6��N�T���F���d;���k�#�ZBH��{��H�X-}�$��;�"��"���g��I�|/MG�k�N��u��߄<i��T_e��s�n�(`
�VA���R���v��p'������~.#�1_pydn.��Q{Y��D5�ZR�#�.Wt�+�*����I��SJ�'�E�f#���� ������t���Ia��W��Ӻe��|��dl;�=�Ѣ�����	tZ��?J����:��18������30d��;;�\�ݶG@�8�	e_4���QS;>
���諗�/B�BM������'��v�Hm(; ����j*]�׎؈*^GhN��!*���S9���n�ﰪ����B�_�f�f�`�;E�  ))��8+�;P����K��l�"�.�c곖vXHc��L{��St�Jxom���Esa#d�%Nf�_%�_�O�ȶV����뇒���'���׿�}L��@���e�+��+G�~��7����/�h\Bτ3o���dY�0�:�%����, ��{Y�n�v��S�d�FR9�ǫ�m��+v|�2=w���E�R����1��9�DAx�d����	�1�R�x�I���z���Ud ��N�.(���Ӑ6Lp�fs�[��9N(y�i^p��/l/���?���UꀒvI�MiN�{%� �DL;�{hHW�/�g�G�	��W~ϼ��u�N�q����1A�|�+��.�ײb
��a��B|Iy+wG�����mkS]<��W��(%��^�z�&o�������n3)�F���9Фx��W4�Y��J�^
�|B���-�rښ��0�����-���"D��3}1�O��� �:��1!���R����Q���vC�$�z�]_O���!���7<�AX��=#�:զ��j�B«�wK/~/�ܙ=��D���80m�S�9�0_�:��X+ .M���~�������he�?�%�ly��t8*�����U�����I�I��_���!��J�m���9�e�w��ش�E5af��W���!]5,�i��zbF<���ـ�	�s�7P�b��{��̑���>W��ȯ�1}|�[Uk9Å�s�
�ƃX#�{�"�����}�#��JTĊOo3'��	_����Y�u��һ���'�:����Û(�'�:��y-)���C��Ϧ:��LW�"XT9b��;�cϰ��F5�O�y���]c�yǛ����Г�o����ב�s�_d��f�s�U�P0������ci�8�-Y��$D�C`����1����ZsXQ�1������\1��'-���(`�A��E���X��7l'`N��l��r������^'e�Y�i���tx@?�R��E(����]�֌4��)���5v,��~J��k�]Nԑ��m7D�������b����)���h*˽W-'6��m�jk ��ex��5�j�tW����!���7��J�z�Ooo	��=B�\�֞���/���H~�G�o��v=��+����4�b\��O��iW���q�����It�l� �V����M�����q�l �~���y�&
��#1��|�p�?�0�d���*� 9��*���#���F�fB96�C4V��y���m��=�_��~��kկ?<��m�.[|��ʪ�$�F�-�?\_�=x�=Ц��'�l�xp:@&�qq��X����||�T�hF�!�w�=��g1���1|�;�I�����^2B�S#����[�T�ۤ'���	����|�;�є��Y�9<�:gE3��;�]8N~*�f�~�_�䫜Bc��$��.�5q�Q��9Gp��ə4��~6��)�S9qz6B!�{��[�	؄~u���Щ���GD�2%3z�{R��<��w���|�F�[(��S.�[����K��������?�?ޕ8K"?݌~T�m�x�oZ7#�];��굄�'��2�˚#5<����I��y��n����νY�M��'8�D���=fU��$�<��RLd������F���75&�l�J�1�1w
��M�b8�"'G��	�Ċ]���#k"�,������;*6�/��1,׮4���(���"������.�?j���Eq�����@��i?j�!ƒ2#~��i�0�����{�N�r�s��:�E����TGJH�x3�k
c��箔r_�s�ò�H���0Y�����$�:��V+����..F��_���SSO��&t|��!�׍��G�=�2�{��ưk'@�vv���Cpl�K3�	��_��O�6'a_n�pT�RB�e�j��Y��Um�9iT@�K_l�Ö6��� 렾)H�|�ú�&V@���P���-X����g�2f�Z �Z�s7�u�{s��،����Z־ID�����rK�ʊ�r#U�eҦ�~u㈛�g�I �#�M�l�Y������v*6v�G��q�|*<Z(�븋bu��r����sc�Qɍ1�4gފ��օ:���+ߕ�%��`3�+�7\���݀"L�,�X8@� CD��@0w+���K�6������	B7o�RP��3�/=�P��V?������6��o�k�LJ��T-o�v͊[v��%I"]���yg�՜uJy`K�;H��3Yc6¯���(m��w�����՞n��a���T�YS8�:��9hF+��u�]X{?F�H���O��4���F@�[}�
�@��s���7�f�~0��S�-���/�g��(���@i3����pv�iJ��ޗ_�H՞��"����ѭ����$��?u�ES�N�a&��~N��B#TH�٥�{Q^w(q���o^G�Tf-ҚF��B,�/��G�nc�@������g?���n%�\�/�-eO�j=����JY2��!���`�ej��� �+c{ <J�#"h��蠧�oͩ�'�YaTą�{�T�=q4��0!�d:V]���X�n�M���?�&Ng�qD�&$��H�G� zu5�'N��5y+��֍KC��v�O�[�;��
��z	��N�σ��h�w��`�%���[��v�]������ /+5O;�U�"3�C�G���I���n��
6b�kˡ��K2���v�Ip��b*��xB��=M[���%�CR�.���q�T)�,+�4�Yɍ����D��볯��C��&��B`ր���13wOz��KŔ���f��Zk>�x*���v���S��kmy�wӶ�}��8	v���=]ћ礨N��5��㤖��G�1�����7�&��%ٛ��V���(U�Hx�����Yq������R݀� ��F�>�وR�w���E�Sx��ŕ�U_^�;�7�tu�X����|�����F-��[	7U�����(�|�)P�zw�b�R1jB�1�J�7�OH��a�(����1�2�H�,o��Yﳢ�x֑q����0j*��)���
 �&F�)aA�l aO���ņ��)�1�����0�$����򓧁�ͯ��a�4bk+-LsK�b��(��w�U���^u�~��i�U%���93��2z����(5�hz�T����ٽ��&č��Є�ـ���e��)(3���J=�8�MH��	/z�l$�7HT5����,dp��v����}�G�Ay�X^��XX�_�Y�W���*?L����n�cm�+h�u���g��*�ډ0�k����$@Z��:�k�Wv��36�[��X�P�r��	E�v�	�O�^�|�#������ڤ�M���{R}�̻'m��ل�]�9D��MJ�D5��9���aY�#?E8�(d��}�ʖ�>����`ǈ�L�Q�[�:�Cs���\$��HZ΍��:�vJ�yM��Z�����4L�#LK���<��m_��7ω�		مJ���V�}�O�#��e�}�*��Z��ov-O|a����n3{���G�á�cn�l� �M�R���{(]�\:���R���c_ �7B����:���.�$_���%S�P�Ž�~�"�*@���i�Z�����ayts����h�s�,W|v����a�����+W�������;evVw@%x������FS�q��f�iqEX�X��Hx���M����ut�#�븦zHYC٧����AWN����cU�^/��pF��^΀�f��(�ss.���? �>3�{JF8< *�C�qj�G���,;<3�����-��֔��;�E��uyM�Qt3e,wr'~)�`	w�3�b{S�P��|�������ث��xL"������9؂-sB㇅H��C)�Y�j��Z��������m��[�f䇏G�/;Y=&��� ��"p���I�/D�W �j:y�#�i���3 ��ԓ?f��'B8������Es�M~��c� �6R���n��JI��[M�g��@��6/Oh2�=�8�6��K�w�{�>I���ҽACQ���{��]퍐�!��)��p��#���d�A�alU��3׌l^�SJx�[iH�G� \{�u̜��|�P�P�II��]A6��A3�{���,Z����*\����qk� Ĳ�_dhx��2Xeq�ւ�=�����L�c2Y���=�呿_����'��4��g(�������Z}6�C���|1ٜ��0`I]��V��c�;���/L����Ya�e|��"ɓ����uz�YL��+F��R�_r�?p�?�(�/�QC~���50��1�Wz��u����,Ï����=u�ox�b�	u�`u�8�0"��\�W�Ҋ�V��A�=rI��q�����o7���|9x�Ro�Û{�?Dז�P�E��*K��:�A_ţ^�����bT%�G/Q���s�&�-�.{���8�a�eL/�x�P��Bq����ͷ��l�����r��n�7#�=9 ���hS��ľ^�ޒ��S��*З�Z=�v��r�� 8���T
Y�xI��>�F)����luc�a��S��"=��J�s˩?Tw��A�w��Fc�;�t��*���"�/f5��&(P~� �V��r5���i�s�3_�C]��*M�v�(*n��j�S�4��9���g�����u��-B���,q�J!�g�F�S��噀�93��@�Y|`>�+	�CK	4��>4#դ��Wc������_�^-Y�6���"�e�m(7geŖɹ�YB���l?�8���B��m5����U�ُ@�����������6��&"��m�V�����c���M�фP��ó CS����z��nj�������
ꘕT�;�y�m�NT�=׊��� 6��C�9(ľ�zn���nn��t}���w�<�m�ǰ^j��m?f_�'�
�z� -�-�����|ˑ�r���D�IC�#R8~����tȵ]�/�&��z*�'{.���;��(���������a)i�<zVs'	R��}E!��9:�J�����T_v	T��I��x�*9���Ai�ʐr��	�oT���H?�wOOh�����D�#�[�'wvل�ߎ�Fg�Er�ᴈn�ZH��oy)���/�È/�g�?,�(bNAC�P��f�pS�&G����|<K���]a靿wKz?�L�8c��ݎ�������Q;Y`G��x��}��B��\�4�vs��V��u�qERhX �wz9C���9��@n�8��AН������fh���M�&�AF����v�4���{x�x�{F���J��l���X��̬����+@:�Ӣ�� ��j
)au�Sm����ETQh��L�T��������2֥����HF)#셍E�Q��䫱������d��w�TAA�M��zn����᧡��lw��RA[[���n���Д�yC���':�d5�C|�\���4"q��g��o�G@�0�#���@p���T�z�26Q�_�I���� |��:icl�:W��W�K)�b�1G���r����>�k�Z4��a��+b��&��ꋀ�#t��o�!56�y�V%�(w���N�{�E
�)-���;At��,σ�����w5�U2f�<x+��Zfv���ŷ���<��ؚ|џ�Y��=e��&͘{h-Gd����kiL,���z�r^:	h{�{ �T�L�	S���ŶM��V9E4ARG3��O�'�;^hV�=
��|�7"|�
}��u�����R�:|F�o��Xf�ҫ�@ x@�����d��(]��v�%-��k�\HI�8�JQ@|(փ�S��W��SZK�5\��F����2S�^�bݮPjUMx����hp�v{eM���i{�G�]���߽F�m]�0��{�hԯb���̌���Ӕ�g�C|���~���I66]�~�J:T��L��C�ױ�~��^�f�-�(%����?&~�a��Q1��tA�y{R+e�\���I�Q��Fz��/�8�3�_Lp8���b�W�Y���כ�;=��'���ے�`>��g/z{�3�Nz��IZf���vTlsuǄĈ`N���P�%cf� [ʀ�������op��qThȱބ)`+I�h�c�$��lh7���֭��EM����y=㼃�/���H�n����w�(@ؓ�!�>���&w!2���/�"��9_"�:B��
<8c��σ�i��[�Tg�����qW:�v�7$��;u%#۴j؝䵻��;Um=�Mق_98-�G�H�	��� `u����j���rU�X���Ng�P���3ٚ�~�梔*��n��G�֫W�o��vcY������+wމ͊��}q�Q�t̕���_�OEL4�:,�cyN��{%��s�	YO)�1#�r�uw��{M�[GdlV���T�]�˖���m��`*"�$�F>�xܕX�~�E+�0Dsۓ���E�W�|��ÍW'����j���B�>Hf?��)��c&���_���|��D��N���D-��_GE���YU�|EA���,~�ԓ<U�wx�����\B$y��_�\�f���-h��:F�C�R����mb�>�H�s�7EJ}��`������+���!�>�/̠�ѷ�7˲B�	y����oQ��'�->�\�g���2�Uχ[��2�8H��x�)��C�$�X�����x��\���75k���K��5Pt�/Z��	B�m~��\��*ɗ�+�Ryۈ��<E�������+G�(2e�NX��T:���Y��f�
�r]�Kb̨�k��p���V87�����X����q6���(�U�w�'�
�]���yqk���<v[>�a�ʂ�k�W��z��ğ��%y�נ�y-�HN�O��%�^�"���K|�����W�H}{�x*[]� f�r�x�
C�G��� B
��"r�_XXO��M�	I*��8�6]Lp+��'d"��b(�3.�j�冡*0�뵛��A�EP��E?��R�������ͭI��ҳ��X��^������:�����N�}�qӢ���ٳg�~�����$� �.�p���;3�~B�}¥wW��#�	��^\�/���`�_T����
��E������e�ǋ��R�S)���Ԁ�f���[K	��]��/R��߁Q�����0T�{ ������nJ}�k��4<\0��0>��F�xM����|^�>2�g�Ikrs<u3�5i��ҘߓW~^^n?O7�˺�'4�i!zR��y��g�x��F7=�yd��0{/��g\�;�u����2���z�e��ޙ��IU'�b��Xdq>n��I�Y2#KÉx5d��9]®������T��8+N$.`��>��ߚBo9���m�86��S� �L	#&�G����`������ ��bn���^,9�_��U��_�w���!�'�ԭ 	"�E�?�"�]�gv�E�V��*�;�x)�{3Y�����7	�0;Y��:�<� lM��WZ��=�j^mUb�t�x����w��dN�����֚7�|M���[<A�g�&���,qj��i��VS��lw*VTRƞg�$ދ�w&$�g�x�ܺU�����L29j�(8�>~�E��9K��ظ�>����t���כ��v�MG�?�֋c���=���I��'C��T��'���A�W��q�Ԭ4;�Y�n2����~��ht����v+�ݸ�Q��������~p�9��یv�^Yx�^�����L�p!��Oݾ�k�e7��ڟRJ���g�v����?�~�Ƶ9���ʛڙ�K�L|���I��H1���3�Ƨ��E)�v����K,\}@������ɉ�鹴86�AP�2Y�ՠ�\n���K�>U�v��><q�.a��+�g_)y~2���
竫t2Yj3m�sp��r�ٿ�S�R��?�v���h˫����-�\�ok���ߘ�O�i�k��*6_�坸�l�]?¤�*�DO�>����c;;Ox�~}�&iӈ���m6���q��P����l�
Y7�%k��U�P��d��#�X�6e�hQFc�[���R1��̈́���������{~�<8<�罿^��sfLY��������m�Rg�!Fn�"	׸�U��|�z1gda~�o��#��PQ�T`P�������r۟b$��ߒ�=��x\/J�� �� ���A;�6�bw+��zfJ�*�DE7�9�����:D��dޭ����_^��4����\��t���>j��� |u [׽oS">;��s��Ω饕[�h�4-�D����I ���6�n|�N�+n^�\����,���z��C��|���I�̍��{���f8�o�����Ȑ��!��Պ����9�Q�䄹��Yy	 Y%Y�"���7�<�|m:�<�z��U�Ǩ@�˛��G��ɰe�@�ac1Ǌo����ˈ۱�~R *�_w㹋�͎����O>�mJ�����W�JO�m������C0�[-��t�!.�0K���5� ����9�m	�A�J}:v�~�oh�HIS�T9�?j���/[�g�PL�8;[5w���PaEa�x&�0�r�W[���Ս����l��rO���pf�We�}����K%��e����yJL����!���j}y�X�o{@_*�;�կ>���ɇ偰�g�L��7�H���.�tI-��Y��9��+e�C�j$#7�#;��ך��p�������*�}M�|l�_��xK{�'� ��	\\C[����%��݈>Ǝb`�@c0����?��ZF��7ed�0��`���������l��~�� ?S3�GC�A��l ��)���xޤ��!AY�۫#�vw6�*t瞿�\N�����3ǔE�m��3{4)y��Y�Q��Y��/��:Y������(�c2��1�$�l�A�92����f�g��&K�ѻ�kD���|f=CCZ�G�y���+�B���e:���1pG�
o��W���g�;�����7�Z�ф�<�5�p����!�M���*�{3L`x��dCC{má��������� 0<5�K��ZaU��ސ�7K̾)5%�����=���,P1�P�f�a���r0z�-�@ �W�}�X:t�b�Suu��?��	�>��O{�+�(�K��T����M��]����6��@��9vYӐ�m�����$A ��t/c]N_pض��])n����W8������`%�6����=������d�����n]!�u)է콎P�������3���v�5��t��Q��Kb֦8z�}�׻@|'&�䶎ĶVJ1���g�sPuΦ�U�|~s��P@�x��z?�?/}��.���~"��c_4RP��� (�|q�p��Fk𥉟�_�0��ǭv�#�O4��,���N�B�E�W����h��uw�0:�^��Y�1��T0�[d��ŦM@
X��k�a��SU���"��@��%��tn�
������A���G#""�5fD�{��_��CdQ:������
��
� ���ӷwɖ��c���,��D�3����aW�C´^0�02�ӯ�%���ֈE����i�1�O���^�m֜1k6�5X���Q���FQI�2SE)2�$��/�I&�)�9��xE�%�ޤ�;ON��D�̡�(�Ib��%<b�M����������p�`�F�l�{���	���G}'�f��9�E�X�	<��ؖrIc�_���+���m�+S�y�z�sy2{�J��TnΩy�����i�����4��B�HX�$��=�"��g��r߿ �x�,�\Wc���$,���a�Ծ9o&�W�r�%S�/��#.M, ��o-��}�o��Ȑ��j�0��T����<�ҕz���b�(,�� >)j�
��
�}�3��n�L�o��Z��k�<ֺa3�H�fH�2%���Y&��f)P�.�*���DPf�;�wsU��#1��|�؝ۓQ� R&�Us*�7Frv@b��:���6��3"7���H�`k����m���$jƞ }�Έ���?�Z)����#y�iξ�r��}fa ��]elK�ue3c�}�b �]���P/�Ֆ�����Ҋ�{���%0�ii)���}��E��;��9�+W�meXX�z�>p�<b�:q�|q�%v�~%�5s��{���ƙ��[[�#���U�_2�����$���i�$�n~�~64'3�:a3�����M��ʕ���(Y��*9�!/V������_���
�⽕� \ON<�d�� 7��Y/8^�L�n��	�//=�"_ؕ̖��8�R'8��x�Z*=ݙs�_�F�> +G�N�-���N�.v�L�����d���ʓgOk�>���ie����A����?��[
�7����[Y��ٲ����{aN`�d�����)X��f�`�1���]G���'5�&+)�:62a��[o.=�:(xp�[v��^�5Ǡ�l��@�� ���V�����-JB?wn�?{�1�L'�{&:��� ���_�5�p|,D֥9��Ρ�T+�K�[U�|�����hS�"3���������R����B)�5D�#�m1BS��ȎB�������ooH��mX*pQ�N�'\)iϪcd���>ܓk�&X�Z��ַ���%��r�W�傫�~w(Q͜�W�CX�t__�|�Ubbf3��C�����76��T	fK�Ef�`;c�]��Y�e���'1�	��������aw),����})��ks����,"�+��fMg�I}�i1[��ck�`JZ2���1{N���9V�u�:Q&yH�'ih�7��������g���8M���(?,?�*X�0�Bp��4-y�U�ND���D��Ḳ�/nC{L��y�D>DF壆
�������?��em^޷v.�	\5��'S{��^ȓGPز��E:5&��4u³6��=c`����!��9��F�Q�@ "�H��!y��t#��I�=�>��ٵV�hˑ�Yf�{ն�Ͼ���e�?��rPpB-����r�x�3T~�����f,9���W#i�ELU��e4�<hX%?"�p���+/eoަ��BiȣWƋ9콁� �É͖<�ð��{76��2�����$r��ʯn���V���2Y��C�n�kAwj﷗������r\��=�����A�#�c�ж�P�Ơ�"R.����>��v�g�YT�k�2��b�M}me��4����-ibv0F�%������@x�WS���T��俑i��I���Aǎ6f�].;4����o��03���*Q�R�J.ua�G�Zp���lM��n�S�Є�/�Pw��|��;t��b��;"ȉz�9�r;�6�}2*���wS�p�G)'� �㬜xEڪ��݁ߩ��Ho�&T����"�ƭ�!�&f��b |('=��&���1�fZG?�)�,6ӝ`�Ek�J^����1>ah?���I�����Qn�[�䝢a�0�٧��"ߝ�x}8�rl���DW�=|-E�
��?FLhzs\�d I15C>UCڠ���$��F��j�� �:Ϸ|"��4�L�6�E���t]A���:���,.w�('�^D�'�
*R���	�8i��l����)B{�����)��%��9E#�SҠ?���5��Βnf�L�"\��jy�vi��D�H�}؃���x1��C^kZ)�)-�ٱ)T��qtp��I��i���(���Q�*����nAj��VZ��-���������;�l���	��V� �!��,>����pr�� �^˦�� �yY�)���!����@�{����y�0�P���]��g��D�b��/��/�7�g-�,�F�;#�1�����B4�ԙAv1�5*=ƶ�a���CTN��b″$��6��G{�|2N���f�I����TY���P��E?��{�=Q�@��q��O��{��֥h@�!�>��Eq�s��'eɈ��d��uW����)Zfd�/���V:tFEqZCǙ̡}�_m�%9���H����Y�6���N
"�:O��[|�����op�
�� 8p#��>zn�	q���,�����������u+���-�P�T1�M���i��������[_���lĈ���	��]B	��&LGRj�*ޓ5��r]�0Z60h�<WN�k;8�o�\��{%�擛���c���Y��	a֝:�(���烣P=]���5kky�.CO�3+��C~�`�ƃ�X����������	�2�x�!"nG����k]�!�$-=�� �Q�Jy�X�V*
Ol[�/��*�4�-tp#͔�%���@(-5�����ʎ3:�"CJ����䵛�bN�3�Q"�9�#��얇� �����4�3�fVX9�6x��䨣�Ȗ+���S�u&[�\��c�+��ii|�;���-E_%��4
��Q5��r���C�����c�28Jr�X]ѷ�̖���Ё��ax�
6(K{��
�KT���Щ�܃�����\�~���HwV��U�0�tt��""�É���:�9M@k�:��q��sj���_D�F��cF����ǘʹj� <{h�����7�" �q4r�[��������5p݅P��Ҡ����_�"��k�,�	h�t�P�=���C�"$Qr8u����0#Y.Z�x�]p������TY/=���|�"
H����?�=N���?�Y.��f4m�T-0�i����ᇼ�9"N#L�b�D�p?��t_?��6ϣ�K�����44JV$C������a�(�� ��/�cm�_�p˗�7���r�����Y�y[M
,�i�����{�Bo�;��d:_������9C�a��DIڣ�d2I�"㔁�Av��9�*G�i�i0*Ù���y��G�Eg]@� �t(1g���G��	m�P��n���K�nبP�:���Gi����DR�Knp�f���>��}`��1�H?�^����R�I=vB	�7V������@�
l	�O#��Q���A��O��=�����qi�����^S-�)�d��S1V78V��������T/�2�l��(�s��d�
5G�O_�rr��<K�iC���S����gi�ڵ����"�W+��� +����lt�#��
����;�����8&'�O�\v�B&[��hs�k��I9�;��op���e��GR��bxAjolث��↼I�^�Y:X�Х-�Y��'=����&�C���~��*����a�v��B�o�-0��L=E^c����"�C�$��I��r區��d'� Q?�)��n�v������8�<,���*��� @���KF73�+fv��y7����P���E׷�͑)��b�1�&����a�0B�FJ#�}ۨr�a�8� pX�����em�.���[#��e)?��MbGO�&|!܏q���m�M3l��i��O=U¢��`9�����
պ"2V�a��Ӿ�?�c��Lb%�&�3,`;8,�A�\1�Z1<��s�*��><bo���km���o9��7wEU�=B'�g�.6Yt?g�@�u�r��������~y����ʭR��bթ&�u�z�rR!�8@{��/C��n����|�Fs�v&��wƝ�/�H��N��U`Y�,_��%|�"o̝���D��z�y��Z P�\�^}�5���5�=Z�0��S*���',�A��z51U|]��O��,��>W�<}U�j@h��l^�"���l��Z����U��M�k���B�.&:4�_�м#\%���곘N3�������T��]O�e���h�0h}�;���H���'@���{��\�-�������~o�t!Z"�����kM�n}[�a�����c�䓷�$@����f��BX�,�/߯��r)����u�h�E��6�ԿڡD�|t=�AOx��*Kt�ٲ�T$ԯ���r;���a�V�{���J��kx�9�}�	��^���8���c���7�����]���IO3�@��e�M��+N���PK   ƮCY5��<O  g  /   images/4c6ee15b-826a-4754-a49c-440dc66ff58a.png�x	8�m��P!B�a�0ƾck�l��Nf�1ƈ��O����:�}�,3���'"#K��NQ�o=�|��������������w�׹]�u�w2�ڌ�[��D�-��8��ᄧxh�0��	��H�ۙ�Q�do���Lup�9� �������S�@)5���MwT�]�(vdD�?�\�	��]��u��K[���mT�
+G�yK}��*��~,�[��>�_�5��R��-]�[�Gգ�/Q�y���_��{>6�;g^bɾU�J���P���H��d+��Vfɮi�JÌ�x�>�?�UPUo*!>'�Y;]ʓt�m�ġ3�-b㺔�Ur��c���sX���^ς�cR	�'�&�q��M����_M�m�<`�S�|g�?N���	�V�{l�Z}.,���t�*�O��8���!;����EyZ��w�	")�~x|83纀ǵw����摧+�9˛
�h)Gbf4�'�I�Z3�����/r[C��k�.-��~�����2p�d��43����G~�x~r-:�@�󧨏�	�P��EY7⅟�'��65Z��ت~wj��C�bS�Jiw�0�I7R��n�}�Z}R"��Q������pT�^N�aBX��l_t�FD]Ь�#���v�c7�����w	`�r������q�
U	Jq��-*>�Do	^w�uk��[�^��{�U'�M�?/R#��J��[�bŅ�^�1�Z�G��w�Q5_�~N���g��~�F;�1x��䌞����jv�9&#:u�Գ�j��*���;�o�qk���^}����-}�P�#��o��f���)|�-���X������gs~�A�b$�I���[/�_H,�[���o��~k�����Y�ϴ2kφ�7�C֩�ʕ���:�&��c?ښ^GwD���nuc��ۙ7��^)@*Ƚm�wY�u,R$�`=�S&���i?aI�����m=T���qy���Y5�)R �GH�yIM�l�nVrdKެf_��rp@
�q\l��l$xY���M��C��ې�);�~{]{���>#����*�}�D����k4���-����p�Eo���}M��l�Ǥ҃_Y^�Od�\��̏�\]�Qm��(��n�{�l�8��4q��y8���;8G�h/'0k�[%�����[�[k�P��������hMK7�el���7ܮ �Sc٨Q=��.ubo�I� �Gp�fe������g+K����%{��H��K� ,�Ë���=qx�?2��������U�	��dD �>��A���B��zap@ 	G� ������a�O�p�}���B(D�h�v�B�O�q`-%����2XKG�S�[����VUVU����T4��*pU������z�퐦�fz�� ��BCC�BՔȁx����LY��
Рp�G�?H��$.�+�@!���;}Or0��K!x��\��_�|���T��a���0�����¿G�y���7. 8��IX/�G��S� ���� 2��C�oD���WM����.$��� �I�?����8�.��3	Ԕ��w�?A&₂ W# *������ 6/s
.@P<(?!�� 6�@�/��q;3����	���7�Q�0��3� �築T������,m���'q��2�+�jPU5��\C�����WV�jE����-T���OP������z��Ɂ$������!�8ΏLHQ�G�9�����# �� �S++�����g�D@ ������izzji�@�pZZPuu�T�ӄj�p���**j��G���w���x��p<?��x��������N�(���_K�w�כ�35�^eI�G�E$����k|���?��/Xٛ��3�6�.q�����)���Yyx�w(��������
�� s`�e�_���K��M��O��t�.�8@t P���Z���̑F�0��<�$��C/e�I������q���H`J9]vYX�r�b'��{v�]A�F�$K���vr���1��<@��loM?��@�����������⑻�6_lq}#�>Z�9�ݴ��`�V	N�Ɉ�O��G5m~it��!�H���mL\

y�F�5bmE�~l�q*%m���ɤ���y��+�Z7�Lo��:�8X�5���E�rA_1��ML�[�u���9��o����¶�Qff�);���=�F�u����t��.��2L9�����G��=>}}+B�aqt�}	�6���7�b����g����Gغ�O3���7C�嶷���WҮnWK�Q�a�_�EO��.�o�i�&V�b���617�=}�������fi��u�{��o�,���0�{������(?	_}��ڻ��E6��v`�����������?�WV�����l�i�؆�>���+�-���{u�%�)���PuJ�$w;"�#�2�S8��������(�Z�@L�.8o�����o�*����ϯ�'�\@����{=Ș8ܷ��7��-�%��+����e8N�=rfZm���X9�uƥd*	��5���g���r��A�?��~l��$x�w��}&�����6��>W�zw��C,W�-TTWy��v92cw��;d����h����`�l����.x�J�)�ą���{e��(�H�MO����[��� �����99:�[���Gx�x,�y������ثu<2u#ꢧ�ԏu �I�\���|�&6&�&����ۧϿ{ZY��.�װ2��#�ĩ�Ds[y�6#�UO�G�v�t����{�y�h�BM*[W/�R(�x �p��K�w�
�h��Qh{{M��ZX6���]W+>W�s�[Y��5�	F�Nf?֜!���vk��F�_�̬��j��gU����
�Ǉ%+<<��EQ�i�M��b6>�L���zf�J-�����.#�j�_�ē��j�H��cIl´��d��Ne�H
��0�n-�������p��8Ց�!�E�WK��Ns�Wg�X�����DҔPHh���Ř7�l�2��`�L�K�L֍�2ѝ"�5t��6�X��(w��c��{���]B:$sY,OU�j�]^���3y��8��:Qa�&f��7�3ya��
ZV��t��I�aw�,������C/"Jrh$O��i-�M�[ �sZ����;�%rt^ߢ/g�hȯ��P����1h�#*RI���h��n�Eq�mE�]���q� �p�-:���i��ET�5�}��2��r�:��COm"���v����'-��4���yQ1���JR�a�!�L.�sֽ�/Q�%:�6����X���5�|M�J�c��8����J�W�+9�^ɹ�B�-���h�H���HΥ�����y�K4�)SR����OR2�G�:�H��W��)�={֓v�2y!.���b�s�Z���������jz�BVإi_�)"�`h[�^�]�ɮG��Lh���4nꚞ@�'I�Y���Ǵ�w���<���r�#���󹤆&�(�L.�vE ��1�H�k��#04��_���z�dJv?B��j��%�{�����8��v78���⨮fm2m5����<����s<;��l!so�`�\`���K�Nz�q�f<I��	���[Q�c�F�m��@�GoY��'k��R'�u�h	�i�(]|?[Yux��M�SE��]��3�\	����d�Cb`�(�G�����yRv�|��|���X��0@i��o]0V� �=�hw:�E�B�C ���V�Ёt�p.˰�� _�e�i1�_-k�S2q&�o�1��tD�r�9����1`�H�/��_0Yc�ka������M�Gm!�ed���tZ'����`�DQq�����n�L�+U ��)d3Ʈ����B Q�5ya�!�F������v��Bg0$C��/�0�r�C�)Oi���`t��bݫCϞ������<I=(C�NUb�9|%�T��
f��9��MZ>���[�"�4��"{��/�b >ጅjGL�һ�,�Y�$D��[�z���|�B�x�,O$F�UӏE��A�"3�+��Lӯ9:E�V*����Є6ߛ4��.�ٌ�rE�C�yz�М��!�ʁ��Y��D�T,&ϸe�q�׿���
H�����@~5ٕ����T֮�G�lU�`�<C�W��tm����V��ɪ}�#�3�hҺ*&T�m��e�V�1
S -T9�ϗa�;M���W5x%�@uFʬ�K5};���~�N�(M�ƥ[�>ټ]w��Zʗ�0�gw��sq`n�t2Ӥ��Ͼ�,#��ԓ���nQ�С��{���
��(u�@�d�!Q��ߦܙ��=gS���z@R�޲�����KjM8�0X@?�<	��;��)�r����j.k���y�Ȳz�/���?^�&U�Z���e|��/�7���0Ԁ-2m���}��*�XS��Ih9s��<H�F��'y�E��ߦI�p�P�CA�l����q�Iwq�^Mʙ ��a�+���5�"�KI�����ѻK5��br��M���&U��y�����Pp�F��|��ٟ�qɐ���q�C�I���D�� �a�ާ���TdD�˩�om:�I���s5f�u�����S�{��I�G�œU�D��b6�#}�Vv(���R˄G�b�#���O&''��L]�||��}'�8&�d�����r���I('��mkÑ���O7�\�-l߅�_��j,�?�1<�FI�o:h�>z��b	5_7Tihd$���3��ɰWv�%̮̭{WK�2Tf�!}���]"9��98�Ԙ�ö��o���ų�۲	��� ��/�y"��f�狥�?����p#Ѷ��.y�>>����?���ߵf+�1��)mؿ0�б'0�z���O��M�R��D�ǥ�hE��G��i�"6�Vk��RRInr��,є5-8�[3����;'�2��M☐�p�F���^�A>q�J�a̙K��U��\(̣�?�>�}~��0�����{}D�xaěw�'��s�P?�|k��h�K��&��B�]�d�ƈ<d����,�`Ij�xe;5e�����w �$.��?�'�}��:�]#a������P�Fq��Pn��6	�%���fw)�<4GM�Pl��а��q����P��Ư��/�� ����b�}�B4-o�@����M��N�G	�[+C�W�'���w�Z�,ߒ�O ��_�}>(����¤�;�sGlOo�Ŏ��,-�Y4�/�"�3fa��b����%���,�՚�!㦓��b��c,o��۩��f�.�+9B���H��J����b!�מx﯎N��[��ix���r��y_����Sk����GIm�[wt܍���`o���L&9�yґ��*����n��'$�?�I�i`�T�#��j�j�5)o*)/�h.h�H|�?����}%��qd{ f�,����E����f����om6��ρh����>�G��v-܊hc��8L�&_�2~��-���u�5Ht�LZ�
x&��L:(�}r�HXJ��>�*�ez��ο�"�������wl�7���$��e�]��bb��bF��uG,|&�ag�X��C�5����wH��vH�,�;�w���ZCy̨����|�㓎U����%r�j��T]_�J�U�|s&r����	ZJ����[��7F�a�jw��W��1�����8׻�~V��GO��Xs�Yǌ�}�V�ߒe����� .�~��dm�q��j���C�CufM�<C���s��}��j9������u{����E6�3�G��m�w�BTz��6>�_޽6�c��P�Hw�.�9#kR��/���9�B�2C�_��R�|6b��j������x�8�Ն��B;���)�}�o;/ږ��zA�4r�e�c�zA��=^���H�c�z���K�@�.��Vy�5�`���F(��Ċ�d��/m,����=f��_`�6��z������ҍE�ݬNf"�������b��ɘn��w�����:c�i}�4�\h��h��vp�qf��V��X�������]�G@����q)�������e��9&�Z-�rLxC�����k�&Ә�5x�t�~�'>���j���-ᯉg�bI���}'��K4�r
��˦�$�������Ys]�m����0�y��%o�h��LMMM�-��=�R��k�}(���Sf�R�JϳU�4-Ϝi"�t�7D�Ϗ�O^}'UG���F��\?��%��?\3������h-}t0�dʈb{�j��tpuCC�jfwy���י����1�*q�ej�2K-#�Z���x����8;�ݰ��q��fＢl�L/�P	�j����l*�Gf�`t#������qp<� ����E�<�zg�Bk��[܃�?��&��{�g��?PK   �v�X�}��k �) /   images/5b84a191-11d0-42fc-8d11-d4f69521b0c4.png��y8����F����Q�%�آ�B�){�ed_Jj��ƞe�Dv���lM�})�cKx�>��s=>�+W�1�9��~��9gD��i��碇 �ԭ�C�Z _�t4���7�'=n�yC�:����y�z��9�S�]w{��C/;���W⑛���C;	w/��e�n�B��/�τ�Fm��=��0�K�n�Oy�3�L�'D�5�A��if�������Cg�Z�o�܇�}-,���Ky��Д�L��R�:&>��U����_u�}�$�An��Qj|;�	X���>S��,��6����Te����J�����_���x�
�*D�o�r�:�,�ܰ����%�&��a�l���ީ���!l��+T�&����^�y��w?>o���{ۈ�������_^\8V�R��@�{`�O�iY
��.��n�R#s�S�R�TO�066V�uG��P^F?p�=�������s��oX��?73K�̋��pQ`�ϊxI��	�ĩv4�4\5F�v��S=����;7f�Nw>��C٫�7f�(��,$ܥy�N�(�Aw����W�/݅����ؑ�<�9E>*0,����`�N�7�|���������~�|�,Yf$�&�+ƺYej�kub�7�g�H�jQBP�p�^������~�Ɨ4O�s2����]E2FF[���M_P/���Q��ԃ*�p޺��9.n�T��DNg:�#�p�X�M�-A�jA�Fݑ[A�|r����:����njl<��5��7�I�zrȧ���QU��Xm9V�J���_�#�ϖ/��"�� N1<����#��AƩ}�y��3��t�J%Q��:��Z;���)r(S���1�Z�)��H��p�I��lS�V��ĕ�����o��4���i���t���T�ܘ�E����-�z6f�.c���J�����>d���ͪ�L(��A��:�1�4&k.��������,
��L\4"��,--O'�O9�F�`�)����'�������Fr+�Fc�ti�"�U
�w�z&�MPM+ԜN�2yc৚����ۿ���r8�6��Ӫ�1B~��E.�H��-~"�J �͔�~��I��<}n6`�'B�'�֧�&3f�4R��e�w�V8��4յ�z�G�F��ttIFw���y�#����7'��0�kȥ:W4E^J���Ȗ�Yw�����6\���5������}��]f,f7��9ʥwAavfFW��af�
�_]ڀ��A����s�ܶ�����w��v��V��~�3�GW��4������R��"OAev�~���w��"�k�)t�����&D�f_0�m\��1'�Օ,걌�`����?���Mؕ[��@�-���៌�#J��N�s6�QUl���Ta�U�Z���wEv����h�|]{!.� ^<�ѴB	�xk�{Q1�NE����P�YA����F�k|��fe�;x��"s9������ب�?�3��7��as�f�I���3�������~+m{���.5����7hJ��������3,��D(�+\�`^#���Q���2t�lC>YҼ�`���&�W��_��7�?������U����)\(+͐�%�Bȭ$I�V����Sw肃�7JN�}1���"�Gö3�U(?�ʕ{�%������yB��77�3������0��vT�c�[¬X�(שmQx>��I�A��Y:�bH�մ�����(f"ҡ�f�vz���B�> ���2|||ο���~2)�KU1i"��f�R���BT��a�;�_�'~��g�5�\��(��RMX�V��Țd�2I l��r˯�����ܙ����"�����A��nH\����u�KQ�P��mkE�ZV��ң�j��ݠ����>k����2㒜��q��?)��|[�G���Oy�`�xfD���pASj�L�����pz�.M�����;�M�sZߠ����rL�2�.gДV�����g#�Ug(�3B�MЂ%�S�6�~���fRN��(�����.Z2��o�~�j�FX�=��3)�t��
c���"�)���w�*A���Nk[�H�w�����B����&lH�=�Uq��ow��m��p�+��C��e��q�	��GZ�M����_#�m��Q�_����<�:�l�r�	
~���]#��䦚�:!�ԌX�`�����Ӧ���`�T�x��G�d������2��������b�U>ĩ�\9Ac,`�0������ؽl�$�tW���4o��N��gi_�=A�o�
ã";	�4���|^ȟ�1�t���6�@�np-��|<j�5޼�}�#8���XX Ÿ ��X���.��=o/�z�%�lm��2�!NOV�:Z�"�8*�JU����;I���L�� ��n$��kT�,O�J��Q���T��V�����0x���ue�iݝ����c��u��X9��j�:⦗�V�R��b: �G�r�"^�W�ELg����([�����i��	b�
�q�|�
�-�8o�����/�C�io��p�P���VP�b��#�����Zof�T�6p-��||�y;(ˠ)yވ�	h�t�{�,#�DaZ�v�a��*��G��6CD_g�Uj~��#����a8g�.�x�P�?����z|�FΪ�n,������^�37T�^@�+���=I����0,��~k���=���>��|��x���	��(��^|^k��.�S��"S�M��#�OU���٠��?(�ܘі}O��Z��J����q�)q�����Qމ���?�bO�X���W<��ty�AW1��;�%2k;��6(�+�C�ņ�ʹղD���{�xu�P<��.�WZ �gM��Cnƽ$j�'h���;��^e��C>jNp'X�PV��Pui��<Z)i���Q�Ş�U�x
���`1�?�B]��=�o�<% �/Z�M�\M��VzaqQ�7\�
��͌ݰ��q�^*��*!h�܏w53!t����gE�uՎ:����*��n��${��k�}���d��|�	�(��ˬ;o���me���SB͒",$�f���
����r����e���^�`Ir̴
��i},4=�L����ּ�ؑ:��J*(�z#�ht�2T��hń�<$������ ��j�|�/�-��]#�ڋ���{�"�~E���_�R�+1 ��@�닸PU���t�v��e,�����&�rҦ�ZsN>��X�U
Ў	s^�A����}�%%֊;S�e`�����Y>GuKA՜#�?��ϱ��=�wi%X���B���1��v
7���!�2Bp�}L�\B�u��8��Z����޹$�ud?G���F�����]�Q=vf��5OVn��I)+�/ն�X���� !n� �?� ��{v#5�qI(��q�g��/?_�/r��ե$�/U������7?T����E����A��FT�[�#������H^΃}��j��)�"#�{J���X���l빵�݌cH���,��Ԥ�&]JJ��m9\G<�n��R#�#ԏ���r�b��ݪi�mt�����":Q��8��T��(s*����j�ϯn 4eu�c䓀�8��۸���R��+(�O�ǈ�a�g�UX�.��u��\jF����h�m�z�zY�e.͏�<��O��Y@-Q��''��p�5XHm�����ױ�9�'!2t{�E5����KS�	׹�K�Px���M�'�4�sId^[�֢��B�,f���ZG����ې8�A���3n�WdgƼ�z��V����Th��3#���0Vw��f�T/Lh.�x�*�\��<���(�.<��>9祸���x�t�g���	��gvf++Low��}����⭊���S������t9���&����!���JP X;hV�x��	݆Vy
Q�� C/�����u�o���.Yb0�"�ѭ׭O�ӕii�(����D��e�;�\}<�� �x	*�g�>E�Ʀq���ד[A��6F�i�}�3G�B�']������������iL����tx���yy
�6�g3�Ee�� u�[6{�T����O���x��f�b��|X.Q�Uu�G�ǿɸ����9oĥn��^�6�?�3Owtb��n%^�@,���.Ht��;is� iTB��Ag�CVw�Z��lg���ѯG"�?�Ӟ#_ˊ�n)3^����`r=��(R=�,��S��2'�y�u���e���2�&m#?>����ا-�>�L��Z�DN_�k^S��~`ی�NQ雷W-��I�	٘��2�΋�cA�:K�ݖҧ���VE�Ƃ��T^���.y_Y���f]����%?�X]B�}C�΅��`e��B8-�k�=ܠM���gB>��� Q��rK��+J,K�m>W>�8��T�)��\�J�J:rxk��B���$��^!��|�`=Ǟ`�]Ti%MMNL��v�V_@����5�>���1���0�)sn�E�xY��
��s��n����*��4�y��|�<FO0}��r����;�9��Qa*~�iΒ=pL�n��)1���3��t�GIҚ�8:O*o��Lk4���^���x5��õ�s2��] Ԝ�s���7xu��ũ�kq���i@>Vq/�gnzz���_�s����ԫ�.�������6ᕈ	�
�6����F��Ͻ���;I���C4 t]�?(���z�l�IS���5�/������eɵr��Oy�5lBqJ�l-R[�n��D�7���� a/{N\9��J�v�-��i���'�m�,������0f1���XH|��@��*�vc�QiBM��˗<��|g�k��W!�d����==hZ���r����F�8Q]�����nt�����3
e���Fkl\?�.��X��VdKv|L�8���w����3��|&"�/����2U��Ɩ��1di�H>�7ML�gU�=ި0 ���g�P�^��E[չ�X.U���a�f�?ux��摁�r�b*�z�����%���'Ԙg��f~b!�ʧ,u7�2��d�9X$�����Q��>�W,��<�Ö@e4�f��R$�WO�*���t�W��f�ɍ�h)E;aOjL��@L�������+Ulȉ����%迁%�Ƨ6doLQz4O��M�@�SL�k����4�l�b���1�U�ҍ�c�w?�*�WS���d���ҽ>}&V3ϵ����j���i����|,�괣jN6��ٗ��������ޣ��С`���Yý��zdT�솁ԉ�.l U��|*�l���o�;�C��R�XM�\�{?T��`%���#.�D�;���*�ܓCp�����T1�]�:םV��׏�o�Hվ�p{�{���<�w�F�z�|i�p��y
?@�3��n%�M�K$�b�s����-Gm�ou��,��DG?V����-�[����������o�J�/�1ݥ�s36ue�qL��i���ɔ��n�+�*@L�j�$\��z��Z6X�w�[u�҅b��\���e�%��{��=q��X��À�j	j�F����dz��y�DX�������BR�TzMW="nX�PXb6 �	�/� �A��.Ӡ�����N$�c��Cl�B��ܔ�Y�F�V444u)L�?�T�c½�tΧ=/@�b��[C]��@enmog���O�&"Y��\��+ٻ�z`b���V�.�M__2^��V=��! �"���9��ŕ�ͯ�Ҟ������F�ٷ#�^
h
��[����O��FP+g�:�#�{?TP��.]ʓ�W���hf'=4��R�B��2�Ϋ�B@iY�Xp&}�I���� &X"�2ż�����
���:y��j�ʂkM��q����GZB�o����cc��Sd���p�&h�;$��˝�~�1hw}~����&̫k��D�~s�gۗ�m�Q�+��N���Juw6K��>��R�oŏ�N����o����V%[I�@����=�G�M#4r������{�yk^���8�%Q,��wd��7(w��xU��⚦W(���c���\zN����V�x=�HU�� P�FOR�+H��}��������`��qs �bʢ�:"l�Gw��A���E�r`jI�CF�g�lS4r�O'�S�@a��=6g�s-���a����30Jd��@��J�"�!��
�����Ǐe�/��m�e���d��������jԚ���pf����˗4���/��+�B�Ict�p��}�����Qv�_��-���h<q3ڡ��U��/��愨��x�g㾮������RԃY��*��Hͩ�)-ᚑ])5�׷���p�?�����y��j���F��H~ܼB_T*�	���*ŗ���uNt�o� J=�����2�uP�G�����ǈ�l���L�$���{���x���~J���C�jYŬG��f��ć�"s'�p1�[���n�$;KK����V�ik���X(�t���c冉#0&m|���eߌz�>0(�w7��+��),���N:5t��#�}����(;�Ҽ�y
әƕ
���s����飋�r���;�0�����b\�s)L�D�C��E���bV������qm��7v5#�T���b�Z��i�*�Ӭ�!-6��5�<{��3/�<	�(����^j�9#뚨��0
E4,�n��Y�}�����wK��]F��W.]���p��4���,�{�o%�s���@�>2UO��e��+n(�f��T�Z�Rc����I�]q�~q6zf�����߻�m{^���pOg��f������ݾ.--m��d�і,��<&��ج�����j����/�O�1e%%b,6����r��R�[}P��@Gu�Y�3�����I�:*os�V�Cb�;G8u������1:_l���H�#��~�UQ�ߏ����Z��ڤ;��y��`N�7q�tU6>�V:5N��E������ 9��v����k��/
����2�E�Z�g4�Gs5����h|,�\��T�'p�dnoi}�˵S̲M��a���	��KA{�r�K�
�sa��ݻ߿�w9�'!$d�3#d勵��ۑ�[6<�b��\���9����oI�����n��[����<b���de��ן�{<KUl�d�l%���[A�8�:�;������%��e�"���2uy��㼩�����Q�*ZJ�EO6O�3�vR����F��˗�cK� �k�� �rrqI7���Uav.�Y�y|R-�ш[�����I�<����A��S��By`0�>4b�+���������8�5$"�Nk�l��C(���5�hQM5-��ϵw�:��E��쎣s`U�]�z�O�:ɛ-|�R�/�pC-�cu�J:/R�3
���Y����vf�MW����VS���XM��`X����!��<%���SZ���p]ɼ��g�B�"j���o�ì��YJV�m��g8��m���bh�ޏ8��Qe���
������3�'����G󩧙��>n4�ț��8-�?2a�θ�S�TcU�\��&r��J�19�o����IK[���� �;�ב{#�mK�D��z�??���tH#hCT�,*o�s!V����:S�q9�/p�������ض7r�:��K��!E��\���(���2/Ĉ�t��d=����5��?����2<;��3
z��$�Lx�&_N�\�k���k`�phV�W���m�����ET6��>��?���^�wp�]ӁKlIv���g&nj�=���AT���[ԟVQQ�t��b����m¶<�R���.O	��{�; #�Gta9@M����ЎT��3����ݍf<r���g9]�-Di���i�)���;ݯ&��tΰ|�^k���]�,5~	�Eyf���k��s��߻OzCGt�M��Y���o�[9C�r(�O�v��F4�E{�2��\�/y:�������K۷� ��I��Ԕ��V�.ˎ�O�3K�q`��r�9��ϛ�������⇪.>�>ZI`m��I�Z��o��3� �97���*N������k���DU���'o�����9��غ!�&���ϟ�r�bQ�KW	M`�v���H���?墽��j��:��;Ŧ�A��␙�+tX����K�S^ck�|\���r���(��P��	s����p��������MĘ��){0��$c��'ĉ�8�y����W�Ĥ�*�Fj\@�1���Sե��1�_*�MV<ܙIV��>����9����P�v�Y�Ι����g���"�j��+�2?��`q���:�
<��]��� 9\�کW;�)���x@��$�D
;��j��6�4u�x�+�P_$c�QV�4�˥'�F�/�������{]�i��~z�W�[�τ�~둦�w���8�u�6`�ϟ����v<�s�`�LX��4�x�fg�B�Iz�[gWS?999���V̈́�\��7�/=��Ɵ���-�G��-��4����[�`�D8��;){�Wye~�:�wvtЫ�d5�S]��2/ێy��8��Ф�����t7���L?�*��[~+I�ux��J��2y�%z!	�Q��(�k6@� <�K��~��n�;F1�bU���M�P�n:��RU�27g�ƽ⦧g�u��_}���A��^9�;�a�T)������f�"p�8t��n^�T)�7���������d���a�).��M{���0th�H�b^,5&�˜��J��w�ZVR�彫jQd�]k �L�C$(�
{����U�npZjw�0Z�Ӝ^g՗���P�Z���3iC|�����\Q��5]�\r���7ᗟ�pIv۟R�����K�����
���o�.}a����|TSuY!��Tc#O`ڦk�똨)�+�,!~/}n��Z|�K1i#�z���H<
+�3�ٽ���5�AS�
}vIvl��������)L�������>�&�+�o�d��:1͂��V�S��'t��Ǎ�wcb�����+0S$D�'dv#:�� -Sa�f�9��B<>��nqe�J�Sg��-_:�C�E6�I,���5D�޺�J>���Wr_�4*�����M������4�-�cu�Ω�K�� l|��^�P��	�;��p*�n�IUj�"���F�9U�v8��DQc`�%%%�g���7m��j�Ds���!
��,�B�>��֙�Pܺ��"鲮�ۨg������R�3^�A��[r��?��!�_� �I�M�S����|�566�@��H�%j��<>~��j�@���X$dc����Px�{�^L7m 
L�p+��������Xn��3�h�յ�������QQ�!�O?���d���|�l��H-d&���'ʔ�-3]�U;�N����<��xqgY�,)ާ�]R��X%��//��=G	q���l�̮������f��0�c~W�^��c�:x�7�����D���ǐ����d�BX�.��nGu���3�=m��&�{��,��P�n��9���<-t��L;`�R����f��`_#��*���L��a�<Fl�~)�9� \���ِPQn��*t����Ǫ2x�XYVf��[H���X)��z�z��+��{�D/�a��C>j�?>��ŒP����$+����5>�<�HJ7��~�%� �Rv Q�i�y����D���'{(�ؔ�.'�7x���]V���%#��V;l[gui	�]#��h+ࠬ�|��K����%��dnU�ɟ���ł(�W��)��@����d���s����T͋�&-��B�0V~S��eC��#Z&��Dۘ�!q_��S]~�%p=K�`�R
��S�Z��é6���D�H+�u�:��|�|l|�b��	��ˣ����Ņ���i�>auU��l �_9��CטF�zgu�tR�/��F�d�Q��`�(F����o����c�HĞ��o�?���΅q��q��u�[68�~JG�I�C���s���f��"x���ɓ'X�i̇��� ��.��9/���]O��:7바;aK����~u�un��a?dv[�U�L�[\�jp�"���~<�JX/ V�a3ˮr��;C!+YLĢ��+���M����H�z~%{�C�o��\��p�5��ؽ��ظd�֙é�������� Ɂ���%B����5'��r�?��mi@ ԉF�7��~�Ka�ʞ[�_TQ��M }�e)�Z�������Uktv{��dK����Ӓ� Ĭ7h5�.�/qX��k]���{k��0���VREe;*IO�=�e�Hp�}Cg����3E(�J���?�"*FZ5[�w�_QV^�P`�'n���)6%S������m%y7�P�&~a�~`�t��Ԯ��Q�`�z]�J9����D�ǐ<���a�2[����8�TK�sC����z�w^�����Qhf����'�M�2/���;o�^���b�t�q�B�F�`�|�l�����Ր�\��_�!��[@J{e0��}�%@g�r0@Մ��/�"2D�Ѭ��o}�W���i��Aa�b��*�O�N���!���yd�F�����R�!�(�����	��D�"L+*�� ߷f$�|z߫6M�5��}wak"Q����M��غ`㿇��6���ed��P�"�}a��L`����Np�A���c��ga_��NP���I��@�=�x�<$��B|�bD*����|�)�7|3�����B��mD�x��_��w�_�|��5��^`A
V�r���1��/��Ԕ>��n���ɷ�v���� �'
�����9�g�6����Ǔc�ݏ�@�l�g�����;<xo���R�QV��#������./=�t��:�
����R��ڬ����m;��-�U��`���?�9�uM���[I�zqY�@�y�4Q��~�_�2�5#TӅ5��{y#�1pM���'Y�_ -]�o�M��:vA��̹�87�����`�2����%>�DF��;���}.r��,_PIE���8: .���~�@��?�t��Ϭ��0�(�%�2�O�������x�)�?I�������~��$!g"�8�rDϙN��I;��ߟ^3�7���K�<����N�'�י��-�b��U�xky�e�jY�7������{`��|_	j��	w�WXN����fQ�m�Ȋ�˲��o��Ќ��@�<n�3.i�[�Q�0��3�[h�}�v{Z��^�~P���6ZP���D�{޿K�p��\��FD	[�c-�k�%s�$ȹ�J�y���*�І�ŧ�/
5�I�q~�Ͷ��97�$��H|1�"��ȯr������2I��5��;[sS�>2v��8��ltG�*k�ѯ1;u��<g'zޟہ��C�����Jx�iI.r����Ϙ�'�͎㓌�ˤ\����T�p|%�!�����V��;&���;1���;VYq��CK �b���#�:%�#����(؅���E�)��`LAM�pV�҈˶�.��x��m��J����+}d�#�຾�R��6Kݵ�������RUtO1���D���t�Rb�n��h�]F��<�!	���ig��6��A�����| C��Un����Ğ���E���J�&%�",���J|��Kc^�D��ž����ه�S��	�U��S���"~���4@����-S{�@�վ�����7�C!P-�{�Ҡ�ә:���b}��� ҇[�-f���}D(��Ű�2Vr{k�W��iУl�u�K���G��-��0X���#C�B������VH��Gm[�:@$��Fſ��:�~���P-�~>*M��eDp�ک���2K	N��TRe�N���g������(,~5���_��+��a�i}�[Z?�������)��A�p"[�P4�]q����%��w�����ױy}] L��<�-�Y��ܷĄ�+��sf��駏�{����U��<�:Z����τ/v1Y����H��8_�I��-�9֞Ț��t�Z�w���ә�_׈����q'��{/tx�6-[�ܿ:�[�$���C�߅��WY���ұ������^��Ew��a�}���S�q��1�B�cۖ�s��������|4����.��*�3N�c���=���h��q8��wQ�}���h��;y��Ѩ}��xϯ5�M�9�]g�����֌�E���R� IzZ��']b��|�_%����D��k��x����I��}�[���3<h#�?D�\�TK� ��H�(���D�35r<^�Ǚ��f"�Y���\ᴺ�x����E]n9�"�+������CwR�μ���1�9v��?�W�	N[gA��AJ�B͂�|��2:���އ~G�qY5XLB���v�)[||��D%���ᲆ��|��{Q�1d_32�2� S=c7���3�C�W$F�����\E\�~���H4ъ��v@L��%[<)k�����$qEߙ���E����� ���Z�[��*}����3�1uK�F2Q;˴��sm�����=����K�K�j�� v�`�ې�`������T�:��pN\Y˜?F���h�1��v��ʲlykkkyff�<e��D���SP��L�M\; ��N�_�3��1�!���s=��y&���X0�2�E������W�N�jbR���:V�J��#�Tb$z�?�T����Jnnn�PW2�9/�۸�u~�``5���������Dv���������V�L�<´�PaJ�F�պ����9y{'Î�x�r ���U6#`�x�;�S	1���fkg�����G��E��Y��M����GONW�1��h�"��oe?����ܝ7����f�}�;	�z����!w���l��S�N�x��V��_g".(Z}Fh�lI�GT����yqB_�M5>aM:w�k��
%^}��ʉ�pyR�.bv�@Fgoo�ѩv�	d}h���h�s�^k�j9�{q�>�Eϋ-�e�}����<�zv�*7�l�P�E��> ��p��}꟥�� aW�mI�q��6����= ����ty������ �����)��p�ٓĈ�"��4�pO�"���+�����)0�d��x����c�/�5ܽW�H8^��ζ1�a��O�h"C�tsj�.���hTE~h?mmp��+��r5E6�;�	����7��� �3��oW$b����X���X�)�#�`gu�����ū�ߴ>U<�t�y��S�c:��F33������܊=<}-�(��T���X+�5/��E\E����/�H$P1V�m�����OG�Z�q�C�VV%":�]�^͢g��ou�]�5`�w=j]j$�(Z5����D�Y;Q���ؽ~h�!�.���sxF���9s&vf���ے��K�,�j0���x�T[�x�fޓ�&_����9��=Օ?? \x��3�Ci�&�`�4�X�. 	m��F�-
��/"�O 6���ޑ%!+��Zd��v
+($L���Xy_�����[:i�B� ��{j��L+P��&
�g��	�=�긯�	�@r����]5<�\��n-8��aP��c�+�A��綵�
�5!���	��f*Z&�b���x`Qޠ㳗������{<�s�5�D;A��<�,����-xn��J���>���YW1 8~�I i�6
h$��8466޿#�zk��~� g�Qg)ͥ4_ҴJձ���R�|}>����a���s���"�]!+%'��[����2�R�L��-��'( �1����"��e�]c6�F�*�D-�z�-Y���tGɤ)�e�!��d����$#�j�k����腫����V"�0�h+n���(/?ono���|)>��܍���M:�o�E^f�W�H� ��p�t�L����2��h�>�%��p���X�I ����|rO��U�Wz�Uڟ�0���M���-�M�����@?�[�c�ASm,� �1���Q��/ɚh\x�G���j;N,a�yЩ�E����]�"���?�4k�CH�2v�x�ۧ��=���DWP�y���:�G�n[�' *�(���"=���������M�{������X����de����Y����5UF�吒!PX`�J_Ҥ��6^,A���T���� !vTT]\ɀ0����&�k+�ӵ[�m�$�`�o��]N�?Oׂ�(z�ͧ�$�2x3�'l��BV�޴����#kȝ�t�I.lT8-3͚ዘ�j@m]����w�G&�^����f�H)Q��J\�]������è��"��E�]:�p.���ooo4�˹Tl$z�wd�"b�y��?��uy��oa�1=x�� w+���'T�#����9�+++�ı�O��lPy6���]�C��@���T苄Z��<Ax{?�C�� �hV��L������|�67����	&�{#���P:&��4����ۏQ�h%��LQX�T�29<��$0f=i�6:��"�4��b����ړ,9Hg�b�.v�R9�8��Q���TTT�BK��Ae-��mꋋ�K�k�8V��O*�����n��[{�a�E`W)b��M�ѷ�f��>��0�X7��_P칗�G��!0���3	/e�k�ב�_1[D�U��h��7�[܏/&�������B�WhJﭡ���-Wȍb�U��fK �/�_2n�0M�uh�k[<���"�zD��; o�6��}�P^q��r?T��������m
xatw �|�8�ə�.%,��9��x���h���`�z�%��n��K�kOmH@��0w%��*����`r�!����Zc�:~�#f%A֤	�$�Gv?R~\vP�X���=���e"������8��nҽ�����Cf��nq�ʼ,w���A0w,��K`%R���T��9�J���*�ד��Y�\G߽����A/�a�M&�Y�dM�Î�{�e��-:��w�z����hƈ $��o�S�P�Y!�6���9f���f���$� $�.}/@9�����k�z���AH����m^�Z�CLQ��h����B��^SP�G<�[���R�����c���-���-q�_6��L��~����14�|������ҋ/�*�gE\u�������`	�(؈9�ťQb���Y3��q�@��:��z�%d?A�/u�by��?|F��g�Z����f�n�5�OBn]M�w�t)�F��GQ����#�2��+a�R����E�����V;P�zŃM�7�oFe�V�%dG{8~�9�Q.�E�����˥�u�KʲsSy��~�շ#®�q�]�ǧ�4Ǹ�@���]���z�m� �%P�h�N������g=�-4E����٣�*(okk��.�FnQB��pO����5J�-������p��uK�G�
}5PЅ�S�Z3���w�o���*0�x��B���	$ ��T�]����g%�<�#2�����OM�z�"~�,v@�S��f�D���Ke�#9�������4ĵ���9<d���WZA$5&�����t,vO�E���<�-xf@`�/��O�3��OG�[�{k�Ѓ��(��� h�3,� -��<m�$�g��bC(��n��o��T7ɏS��]z~Y�n��nsX�ͨ�_�U��{�la�(Wy�.�fٞƠ�:Qh�\�e�`eR�����<=����F{���#�jw*����]d	!��U.�
㟍n,W��SL��6>���Х�4Dtz��H�Z��"4~����y�9�#�:�Wx�S�����a1����k_�8-�1v��!�����.�.�͔�Z��3�n�s��R�KCA�#P�ݑ�����6Ϯ8ު]�Y��%�o*��<+tdG �Qi彙�N<
��^_6n��|���ոY�b��X�[yo�Eؽp	b�
�T���%M��%k���/n"�S��F�2�o��y��k1m������~��ElIvU��w�n�Z��?�o����M�����k�|��#��?Nk��$s��v	Xɸ�����o��q�f�V���N�^U���c�6X vTJO��P4Qȃr"������t��*��z�h�^����q@�M��/+�ՉX�࿯z(GŠ�'�],��޻A��H��� [ƂB_�
�v�	u�����OV����+62�`0�S�+�^����>�B܆Ӑ��5�`���t|�����4����E�N������$�9�6A=�:�k9�~-ǛM<��E5���yn��2�uS�v��}J$��?~�1n�������<���������¦h��Fw[s�>ut��F>EJdlo��j�/�p���Xk�>
S�'���@�F�w�V���/�Q2`0:�R4Qb���{�rf��Z�kP=���T�\�������g��]p�2��'K}�����{�A�1B�u����AǱ�� ������?����3ן#�1�2zܥz���+�7��Sm&����m�y�dNwF�T�B �w���7V�	�[��aԘ��/������me?�.ý���>u6�ױ�l�i��[x
�=�lz��W�P��"�px�/v��(sUY�%`킎
��w�`�����!�v|��.�&B���n�8F����E-�y�(z䁭��T^�L\��9��y��$�*���tpf��L�t(Q����U�[�&r>dhΗ�e���ѯ���M˪����(}I+(Kr�.MJy��I�>�"����Uwz�d�t�ЮR���
]��F&���ƶ����1b�� �q��BPr�N�>E�bzz���ND���`U�k�56#�&�1R����I.���4'�S���C�`������9��������G|�����`$��21���9�e�n�<��%���29Ң:��N��,��|��hs�2����QMm��'t� ��(�4A��KE�)
�k�MP	�"A�(A�H�.Ҥ!ң������v�{o|���O�.k�9ל�������Gw�K*t�A���v�W���
��|��������$6��$���38p@8�Eh'6��Jd��b�k F�l�&_Ek4��Y4�èqq��֞zL�$���1P�]V���g�b��g7�P=�@D��/2s:�$�D����_�)���a�|	ǵ̪ښ�a6梪��;7���]4��e�PGd�X,�G�N����j���,���j
��{=����}�s-�	bUt���&񽙷��O��7����s�ј�cB2EA��ў��7�xPi�I�\l��H��%�=G�������ɗ�o"����z���gx*ls��2�>��[c첯<��f~�()��.�0���aB��L�o|Z�{��j�n>s^9�z��<�d�h)���5}����v�
%P��u�o��o]d�λ�ވci����#�����G��p����?^Y�
�
����Ew%�^7xxt-���S ����XC��g0L��K��C��փXj9c@+��R�f^��ݪq� HR_خ6���ـ�%A��"'~�����3�4��T�dAh��_�9'}��j����ƽ�®�)��/ǔ��>��e��J/5����K�����?�t�"<������"Sq_mm�	�UN�VHUq�V
��R�KkHH�9C�p�s�]Za�����@�Budh����f��bB�0�9�������kc�y�b8tp�+GC����U���k#̑r8�����k�]` ˲�Hz�����4��>`��h+j+��	'�c��6��HK����?*������@�pױ�G�|~"���ڷ����GR����|��j�2�=�J �u�N���>��ɗ�|T��7*3&lZ�ŕ'�}���$J8[ֿ��V L��
���V�R��~V���A-}�4�Я`uTiY~6�,��(�4x��w�v��Mo�����V�u��M��ٓdGǯ�x����ه�f���r�-���5gg�)�A9�;��M��H�!�6�c��S'���ޙ9�zZϒ%�סr١���͆f�c��RW������=S����|}}c��!I*)��߶�M1��Q�N����Ԑ����Z���)yW�$6�g�5U���
��ۙ:�������bM:$�_�ne�a��g����[c#�"G�*F���☣O/�p^)ȼ�����`�һB�򩳴� 7fL@C�H���q{s�n�������沊�ǒ�9 ��`�3��L�mmmi�!��������휌��Z5�hd�d7�����S�$�n���_Wlx�|�����:&e�8��ʊ�&J2�ݖF��?ۘm�K���[>{��$L�h���#�J��-�456!�W/AIӣ	�SS���������-�Bg{|"7/[��/w��a�߱	H�{k���J9%��M�=�������Jm��9Z8���jJ�+�<�!��������%��X�\I~z�t�/%��>8��W��}��Oj��<�)ZE�-�tU�M����j~_���[�K����Y�ق�Xd�$;�q��Vf��T9Yy�f=0��Ywh&���_��q��o�w2���^4�֩����cL4 �g��S�M�<�A��.�d��A�g|�6o;9;gdߺ�tڍ[}�]o=콏����.+�Y�k����d߅��@���N�~m�+��?�D����J^<���\����,3��j�&�[H����.$�:�~m�@�����8���2[��,  RF�!"i�?\�ԛ�PуD"K����vڊq]VzZ��������޿�����Wq�v9�yϲyT�C
�k�vM/��]%c�Rp�e��un�����Ð��6��x�#��y>�p�����s�A�ݙ��[�����|�z�2e&�����M����D�oa�Ծłu��H��lK@�:.�c��P��27��GK��s��z0؛��3�@U��������ʆ�T7߈X��2�b▹d����Bϕ~㕋\P3����'��C��l\��`��4��:�5ũ��ٸ�.�!��Iɻ�Ff�ZU�ę�AM�U�V��@P<N�l+�� z�X��M7�N��{�+�WDH��`�3�Ď�?�S��P(�q��g-�;�����e ��3s&�}bkǑTw��R�����$��1��'>���8�Da�/&B�Id�c�����z���'�D�o���\ή��o��a�Xf��>�x�	��XR"�rb	�c�"�L�g搚vɵ��� �ڕ��s��>e�����S*uqr�y7��$�6Y[mޮ�L�mFBz�G�x�U;	z
?j�33���&�}�,BX����<=i�G'�߈p��A!��D�݀ijj>ґ�F�r�;�����K���8���H&�ȳF��=c�"��9�z߾�0Z�P��_��������@�a.��lG|b-㏃c&�]�������/_z���߼�����qo�.��^�JJ��%$��7�`�#��_X�N(�&�樝���������a��Q7����V����E�(�t�2�}o�c)� � +���f��=�9�f�i2l�&�}q���!�@�g��ÃU�?���f���٣�-��K��`6�f菮M՗Q��bY�n���9��xlV��E��ƽ`ݣ��k����MD�l�QM���M�#{5@u�����z���$��y{�M��tb����ݻ��d�ȯQp�{o�.F�Z�U����'|�w�]�wrH�M�S��\y!����5�M/&�(O+v؎��3��a�2�J�w�tLw&M�<���}�_y�R�9�U#�0cU��?�(�~�.��$j
�:��D<�����R>����&j���Y�(����ey`<:�i���-���p���M�~dT�1��ګ�bi��&�'�Sb�j��3=�s���XI7U��4}j����(�¥=WW��Y��]��QB�uA5�O�@�:×AЋ�XdUBSX�7P�q�K�H1�@ьE�|�Wոdl$�c�.;{8�A���>2����?��x|�������9[��֗2A�e��<���_٭��eKzd:�h-����4��Ǆ5<�~aơ"��r%�F�=�A{��T��Y����e��L�s�(F�+i������<|jt��=�?��4���lh��}?��gYн�.��� ˨W�@g�Q��9�����dG<^��]+99B�S��S*7X��zvW�(oԼ{g���
S��eA�s\�rr�R<ދ�QCF^^�[�j����|8�Ք��=CN�L������!.y�������uhD���W�q-��uZN���i�yY>�-Z��{ޅO��p���O��!!��/�ȸ�d����N	}�j��T�۪֣����ˁ߾�i��S�^����m��ᢥ�[�3'�_ �y:���Xׯ��~��c�S����ӹEE�tuuK��_��e;Ҽ�F��B0Ȭ�O,� F�Q�1cZn�z璗���z!��C�WT�%�o� �=ΖG�XM����L��G�D� �����˨B�̟�<��i?�7����EEW^�\����\��0-��w$*^�nW�=��5��WD�������M.rNkג	H�y"T���)��h<����
�v� w�Gܬ)j�`F�)���<V�!==��[-:ERʆ������
�3����f-�s_4��xK\���-F�y�f�J��������/�J��ā��/�p�+6����s>�{h��J���MV�Q��{��}�������{�-!�X��Q���
��n�G�l[d4�p㿆�W�d��>�(�_�B�����g
>�f��M�qE|�:�YUʜl�
�n�j���z�(��ȟ榍Z���b��mR�gh���Б&lFovv6f��Si�P�ߘÃ��"�(�z������'��W�z���-1�VQ���w/m��h�#��u��zT�׼�b�P��#{?����3(nІM��>��� y�`X�R����Ngyy�E¹�EL�SQ"��F�3��\3��Þ]K9]�I_��)�9�ֲ�U�T-��W=����F����>������Is4�����8g�������N�����Pd���,�2�7K;J�m@�~�K_P�b�,�$�qH��e�;l�������K���Ë>��h4<�Ĺ6a�i6��p���^�A�(x���n��K 	���?��j��U�Lv����aK��&0��.E�߽{� ����S�S�k1�����6qߛB�JY"����1�����/���Y]{�<���r��9��j�VVn�B��(b�d���>�k<��&�_(�$��O3ڋ��as���K��Q�B������ؤ�,I&�}�a�ْN�^��.�1�Qj� |�fN�̡�Ë�Gz0���Q1T3d}��Ro�1, �2J���¥D�3��
�[Fo����'��.�=�����}���#�	j���o��T?m���!=#�ͷ�)��9�Mu+xQ��t����TX�4�oC'��D��SS�¤ի��F��EV~��P):t^ܵCD��I��Dh��%L>�hy+��"�|�]�����(�-eȣ��א�Ͱ������۶&��Ė9��cUU�$"��Ř0��2��ο�g)��L��;xR٣ʱ���lassOK	Dy��/�N�9�%���V�i,"��߿OT
S�"uv�a������8�0-'	W���X��������R��V#}��}�}�g)�ɽ�i�@f�g�)x��:�9|�@C˃x�8:��l߀�1%�9t;�b��a�\"7}��9��k\��@i<�w���y���(��F7�ɄiO�x�w���\p�'_��yF͉҈�D�����%H�,��!!!�Q�4������ k?��oU���_&nz�4�~��Fp�bf�E"�Zb%��������NXr{�,�t���.1t�[9����l�\���wx��R;��)�L���wG��Ή��kꍌm����7K(��\DX^m`[�N���$��&�
9���Bz�������L���R��o������r��7r(Z
)�V� �;���nzv�?�<��D�m\n2
|&��݈e~Y���OT!��N��}1�ț�@�4��Y-!���x��S@�w��6���[�h�W!�6�D)z�dY|�j�
�c�I�K�a�
솜}g����D5PR@�yY}���H��-E���r?�N��o���m����s�w��5H)W�l�8:�B	m@�!�oϜc��y������6|�~`�c(�"�.��}h8
�j���L"�<�ػ�Ū*!`��Zꁒ�A�*���e�a��_�-]����TY��2�Y�yjS��q��ېz[��
gaL ^�j�^�����N�_ՄFy��n�H9Q��3���ǧW�#�:���Ft���K[s� c��c�{�'�r�"��"�F�8Zr�>R����FΫ��tЄ����g�ֵ �r�9��
v
�b�-��S1�;���*�- ]��xlN�/�j�1-u��E���"�6�&�I|B���ʁ�(��J�!~�r�����!��罿�>������|���)U;s�<8�����D�	 �5�L��+�o�l��ީ�<�k�[&R�6&|�T[[[V B'�Ͼ�N���`b>�J����W��D�[D��K5�,��'"O�<����d���G�;������h���E^�E�3���򼇞2-���V	�z`�p�I�[�m���'��J����"CX��U$P4�##2��!���vz��흝�{WaKK:��ͧ��.�:&�����iZ!�2kA<�j��OmvO�?v���>�{���X�͋����:�\b U*�x|S�P����eȻ��]C>&�Z�����t˙j��T�&��Ρ���B�r�|$�r~H��D�cZ��M������>��+W/����E���%C~��%P ����7��E ��ɷ�'��ݭ���QQ`�x �գ�4��bI��!���0�r2c.U�`�Gm:5==�X�HE�;�1�D���&�s(��e��;G��'����R�s��1��I�x��%Gq�L<^8>.���U�b�����yV�rBE&�bq=��m�Ou2���!kI�c�7/���
%m�����e���������;���_��͐�_�"c.�����O
�F��L��c� T��1ܫ���#u-�:	�1�� ����c������Vx��-�W:�XοV�;8�F����E_�t9U��6ߩ�>��jÅ���Y�Db8��k��ݶ��U8hZe;υ�b�Zڀ0�e�h���~P/�����M�%?@U��������:�H$������	?h��;�M�G���,��X��<H�t!=��La�3T~N`Ƅ$�X�� �Yu�`	����|�?���p�;�Ӷ�\�9sβ�߳{�/�>l7t�tcd��i������ʱ�g�3�����s�ݿ�-�<tQ�����F�ЖM�5\����
�X.|@gB\\p�H���AW���kl)� �oOz^S)�4���ؘ �L���	fAk]3�B�r$������50G��Z��`-�>6+r)�rs[�ld6**��Q�x3���[L���b�������_f��B�������.����<tm�F��/���/��
6���.�D^Ax�
S�P̀@��p�]�G+Q8 Rh�\2Ui�� �k�2 ]ﻊ��2����>��r S��;�+R��8pe�t�N>Wj����f�|���k��@�U�Ƹb���7լ�m
��-C	�"�)��dp�2�VA�L,� �б`nR�t�Ԗ������nr��~�HZw��J(�q�Q�5~�^3ȍ>��k�4�XP5˟ ��8�s���AX��RP���s`
�`}���
�,���Sƴޒ�,ZA=��(z�U�C�/lW�|��7KS����5�
;M�n���^ӌS\��&�ן��w��ӄ]���~;
5ebueR/����wB/����<�jS�uC]Óf������1{�R7P_��3-���m����S=����[�n�>�{�����ef�	�6۸��,�K��N��737��}�l�ڂ4�?J�)�����l��m��8��D���e�f�A��`�E@�z~�lj[�N����&�F��I��ALgfkk��ߡg>�b��++Ƙs���@��'�Zq��h6�z�5$�e�7�PXP[?��;���k��24��a���� �g�Z���Ǫ�5��m����5�rs��:z��4�FcpIsd(���_�h�B��n��B�"����ǡE�/����NNeN�V1�(!�p�h�]�m�MF�a��J���,0�ږ�WR��U�I���u*���ׯ�+o2�=������;a�a��񉉁��i��1,��cQD��>��;��7��Q�T�����@`q^?�)=a�X�}�2VY"H.@H@r���X�~�VΖQi�p�,�q��O����ʮr&-{<�����Q�����qvt�\D�b�e��#��9/E��/ �J�����"�>KYd��!�����7���W;�)+.^n��ʺ_R��S�a�MB�Ǩ���k�me�,���d/�^}�_ֳǽuM�'fE��@�?9�w!���
��גO�_��d�}��?��4-���9$�^���S�U�o늋�LL���n�(��O��;[R�F��g[76���W���[j@�Xf�߀��:�\y�{�"����9�}aS�c)�m���Y��Ȓ�4�B����ӧC,P�LB?��9��|j�־n_QAv`��ovh����Q6u�)	�ߝ��v:�t�2JH�wq�d�6�ᣀ��=�R�v�����kFm��O�#������^RJ5��=i:�𼈷�H��&�~Xl�$W��㒣�Ϋ=�{�1��gT��,��%U'��40WW�M��/֞zp�j�Ʒ�W4ؔ3u�e�M� �mW��
����s^�����v���I�w�A��C�;/e����?B��v����w37��ۨ�Q��k�<�͈�y-�9�K�5y��UZ�&�>ִ�,���Xk*n���������i�n:.X"�[yI?�~j�?�2V������I�����B�ӌP��7��X?��ƖI�k���,,,������p|X��?�Y�)��L��xO�aD4����ݡ�����o�0+�t�������uM�p��1�?o+�D>����D2�!��		k��L�M*T;�u#؋}����ey-��;��{��g�(�{�a��'Ȇ=�*�m�1OPO25�r��B
�F�U�������`��^\�ތ�>;��]��|�:���N�a����c�ɿ�� -d���=F	`1��aN�*S�ѳH��ߕ���0:����I�2H\D��K�����Axn�Z�� ���p2>�����n��l���u�[D=~�}5��g��+\�l�����s�f��Q;�@��_$�� }{��u�b��q"5X�����zK��g��K��ig�ʠ�;�le3���HX����ϱ7oހ����2j$nK;;�`�;��cUQ6N��=�s��=U����Enܭ�Jo��6��u��$��x}�e�]E�M��6�6�,-��]׌��p8/�i\4�͈��������m�V����P��������ې/��$������			\�/��2����iү��7^lI�i}�L��|���
lW��\�`�<~��)�0��������K&cZ/y1 ��"��*�][@��<	-�=���
{���Z$�7泌�������k/,/��]'�(����L�臲�P��T_j����
;} _`�Ҷ$I Gfbq�9ja7ES�61�V�;�TV�2��2��`��Y�Ko[���/(� ޓb�1����Qj�żPL���_eU5�z�8��� �]����Ra�H6�%��6�f��7C����h������ߛ!'@�e�d���Et>K+��d��8�k��r񩹾;	�F�h�O�Ro�t��`�0��d�f�r{Lȃ+�tR4n���@���A=
�̻�a]Q���s���q�B. Qn_J.���C-(��ӈ?�r�)��kWR��֯�H����9�C~����ʱ`���Z��d�X���W.�ſ}����oA�����w��aW�Z����{<x�9xx�+ρ���9�ek��W�gn�p�2
m,.�'�*a,@p $ ��k��EGU��9�#�������7�0� �����n������YF=�lZ�q��cU����4�r��F��L�� ��D�5B�|���'��`:>w��\A|��r!b�0S�%G��.�DS��H�Ц��y���ݿ>���Pb$u|�<N�����	`9v?�۾����p9�[ҫ����y	����l�����LI�%خWIGq��[�E��5e7b�=��S�h�F��+�7]x	�����[�{ F~��	ش@����P����a������c�G�^�ڱ�~��	�Y��h��K�������	�5^/=մ>����3�ET7�wo�3���9�/��~��QF,�I|b��Z��:^��&+�:)�����N��nC��D>�k��A�\�3'��Q���"Dߢ���.	j����ئs���ez�_~{���G玜�{�!��Z�h)P����iY�
P+�.�nv�c�w.%�)�k�A�L��kβ�!_����L�j��]���W�@��Y�p��9ći��U��v����QStB�Z
(��E�}b�`L����ҧ͈��U�e��<� ������f�ґ� �&d�|�I R6���1G&��9u-Ϩ->��󪣇)[=S>��0�.�� �(����d�jH১sP�˸�t�?�7�,��)w�\)��$��8\��E�b����ࢇ�s���v(��]G\�ﾌ(Ӹ�\��[�ۺ�ܽi����SWa���͂U�0"�\L�}�3��Ϻr"�tT[	�w��RK�mm���d�����&�4��]��򼒢#Q>:]�/��zV�\8N���cd��}ɍ��_����>�lZF��1k��[��)Gٽ��YC��	t0� `�^�Q]���|��x�0�؇KD����&��R���D��r8�Źܡ\D�����G��B8���|F��<�'��"S),}�@�vSδ��V*4?fhi��pz�:S�cq��2�P�ڲ����:Y�]'���9C�q.{~���PެeT���f?�]
��F��o���5LmfP抑&%h��I9�,#]��}͓�[�ܧ�/��2I��df�o+�Mm6�j����Q�K� ���}��ڙ 0?�{=J�!���'�3��0'�&�.h~��@>"����3q��D����Z�|�C�#�vLz����?�	�cj�<�fg���6|3��QO(ud�)��eߟٍ]D��
��A��������?�(b�{����Q)���������E�ϡ��SZ�?���+�����t�蘦�'�#�!:F�������#�i�m||�h[c�$�B��=�כ�.@�o�0�z���=g;�!e߷D��;�
���d�g7j��~ �P���]5ܛ�\�T�����g5�.�ֹ:�TL>T��3��_v!�@�j�$��E>
��O�݈S�G��I�����;������1j��/��n4��92���v��-�dK ���(UJ������E>��F��$�.f�g��Y�L)�G]���nB}�k|h�����0)c�G����֠f=t��� �mVi�9NHb��(�K'�H�5%x�Vu�Vx�=��e�H�;�µ��)\���E.))�dCF'|�	�Z����-��!'��i�z��ꘙ*��o�<�L 5���O~^/3�����&�!�n���EP������G�����z���1Rem��yAɝ��?.7�YەU���
j8��?a���39b�=z�;s�q���q�eדn)��dAk���m�k���Y뾪��/!f���F��Eۋ���2�^HFçf�w�������T|�:�b r	�����W�����~����)71���F��0����1��v܉��:����00�
C�(�J��Ͻ����cqK�T�br�1�������p��"�h줡�KV����yJ� �ah���������RA;.�[���G�quJ):�� ���"����&nxJ�^��O�U��� �sOZ����t���g�rqqq�|-M��3߾E�y�hS��8%�ͺ��1�,��� 6ñ�к�Xʭ+��J��Ew�kFkEl!�ʀ:��(㸲����Ƭ?�'?S*��_�k��e��J���_'x�wz����u�J�\�]o5��t�����ak��s�߿�9�Dw�@��]ӧ�}��N�L6ۢ.��δE������;]2�?OT��#���--�i�)��̿��5UU�d�uz���r���j�/�>�k�z��K��/�q����I�Byц��_=�`q�~ ��fJ��x�Uzo7�"����v.^%��d�s��Ӟ��`��!T"��-p��P�ܧ�V�uJx#NZm;$l��7��!&�M���3��6��9n�>��-��:��ZJv!I[��0/��8��w�0�Aj@�
�$�	9)�M�Z]XGq:�KXԖ�z\����^���k���V��͐��a{��7�����Ky�ޟ��G\sK��!�AJ�f�h-��X��b{����)���T�6��Q��Ԭ�}7^[��RJKT���M�kkBxΐ�H����y�~f��O$U���ܺ�����[��F�����vv�K�b��v̠Ď���Xd�z(��E����M�X�N�&/!�u@��E���lIBm�~cn�\yA=��xώ���j#��*�B��qp�\|Ύ�;����g��]��
\�R���~k�u�Z1�F�6x�%��l�ڵ�5+�j�/��4����D�m����V�J�sX�#��AE��ϭ����Jm��6$����@��u�p��A?~�|���hI�Pg��lRQ@����&h-��u�T_Jg�c�7o�S,�A,$�ݻK�㈵��xmz�<|7um���$��.r�ߞ��i��N�*5�:	�Re�^Ԁ��w4֞�����ʾ��������N[I�������)���6%��Uy}?Y�]��p8�o���_C25�Hޝ�Lq��"F��ɴ�W��$��2?
��!�jNo�\��G9�T��/v�*sʷ`�v�j���"Ā������ʛ �����A���(�U`.oS]:�ޛ���%*k����B
%�����9�F�b�����������e Lg���С��v�i������'�p���Ҫ��G~U�
CD1������!0]�B�f���(�@����ҳ��A.BwBD�>4�J�1g�Y��YJ��E�"JUڥ{�G�u�v\�g��i`N���̌��olltB����h��7AC� �
�d�n���jN�/�%F�A>jPx�_�>GjI�pR�����˜"p.�M��^u�})��0�j�zh���h��!���ӆ�#�����y !��Pz�!>���`nۨv�7 l�Jl�X�0���>= r}f@y�*wU�!3�4�J�a�F�Z�hg����B�,,��2VI���}vv���%�5�Ϩ��(_)	b��M�?)eSs��RBnjm�QPe��|x��!C����vJPW`)�jp���'�������Q��U 3YI�^]z����Cg�a�J��y"�P��m�6l49]s^��X|h�,�i��-*L1 #�IO�C���R�Y�(Z	0���[��̉VG��L:U��6�+;��F��б�7�=9>J��SJ����m/����at^=���}�{݉z:|���N7c�柒/U�)&Lɗ|J؃�ZV^��%��9�wmH�7J�ii_2`L��բ;״��!u��ͯ!f�/Ϩ�/tM�iZ�\�'���FD8�y |p��i�����{>��tx����Z.C�+]VIc�,.>BK��Ĳc�j?�4p��J5ԵĠ�1ױ���C	TJS.p!�۸�>�/�D�k��bi���� H�IꗬqcB�ˠl� �t$���3*SmQ")��Fw]5t���0;d��
aye�&1� ��R>�&��1m� s��)��ʺ��
�5]�N5+3l�]j(�)��l��1�_��m�hz��&#K�1�8��p]��x ����Ɗ9o���UQ�\��^�`{R��S��l�Ļ��81�3�Z���� ;"t5c�x��{񀒔���R���d��e�'Hu���}�(H!_��p9p�)�@~kh
�U�Zq<�aN��Ca굾`�~r��)Z���d����4�5�yF�Mܡ2}T�"��i�yRx�bx6��0
��	�A���?.c���y#y�����J1�M�߷�ǉ�y�i���PQ��\dr>�������q��*�IՏͺ���t�*0�@,���^��t<�r��
	�;;4?��b>�!��'��B{c?��.8Pe�?~6��B5�aޗ��l>We�0�f���8�HM4�Zc)5���W_�w|tP��sJ.t���)4�O��ɂ^vr	��0���c�1�}���#��F��Ln!�/�C�y�M�F�(�f)��������t��n$\�e�|o���������5�$����m�����bH����r-`;�{��p,�"�o_d'Bi؅��*AA�cp8�@��Evy2���j�-7��)W/�:���̿};�5z���9NtR��43�+(�����,kap�~>&c�Pz6y�~��3�<�k�TR����p�~&�������aD^����n���H��ř;��KW�͑�;�s#���Id�m��؇��bg����C@�N�l=�I�7Q�:G�(�,�Q���A�`�){�#yp
S�M�[,j�+C�!��&Q	��y�1G�ӑ9���7�w�X� '˞��p��#�5<�@�!gK����	�^�an�rt-�2���ć�J��`H}�6�Nb�����h5?Ȥ
y���h�S�g�G����6���P'G���?��\��#��gt���')���򋯰����o��KB�#a�9H��TT�8s��~|��-�6|�5n�X��7�f�>���Q�x��,���e"�����g@��9A=���I�b�r��� ��m��C��,n�����_��۪�+�F��!�N��'��"���Z|�d����Di{H��T����%��F��5[f�)��Z��*G�{L��W�h�8�r)e�� ܮ�NX�+|�#	*�^�}�����$r��x�=?�2��u*�DQa��]]q� [�S�G�{���>_.����HQJ_�0�8�2�`����i� R�Ԋ&H�{���'�.�yL��c�u������7P�"\�͎NN�qYz���*����@ٟ�T��n�+1/el�(Y�B��x�e��ag�@���ʚ�a%������xm �ߔ�	�a��e2�T�m�nx�Pn<���,p�y���[����B�>�uJB&yf�7߂A�k�����W�F*]���(����6�wBNR�PaD��*����fyv�R��9����@�&��������Ε;k'�u�	<Ѩ�F�О%���F�1O_?��JifUg���oll����n�����*8\�_��G#n2��a�WVԻK�=����4� KZ�C}�:?�_�f���j�����23C%t�d��kH%�=J��Ge�퉊`�t�d�	��˟�&!�S�\!3'���g >�o_X@�*�r���8BV�;�B���\�O���+�9M6��&���G��r���a��K�8f~�
���Y�I�@ʇ03m��|�`�'-(jM�`B$	��+���b�/���;�?����1����EE�py�05�]�t�t<y�$nY�_Gj�V�����[��3�^���[E���ć���<�!W	�tD]�0=�_���'Q=:���=^s�象&�v|�Re�Գ��_� �;MC�lI��9:�@o���b��?��K8�|`&0�������xg�vP���Z4V�iK�sթ�o=}|dZ�XtM&T���t��jdC�V"Wl{�A�N�b�h����k�} ��é�[l�����D�0Q/����<�vM�C���,�\E�v�z�65�n������7(��飉���zlO,�ň ۑF��|���)�n�!}�Aӎ�=��H܃&���W�[R��FO
��5t9?�������5�9[x1��/���6�6}c���V�`@!Z�Hԩ'�۞�;�
�����:Z6,;��XW���u$�[�{�(b���1(�x!��'Vܗ�EX�s)F��� �����.OC�p�mǱ�ߗ��L,�@5y�%�E�M�5Y��N��Ζ�������Is�t���+�I,\+�+���1�u��
3O/&w;v�[�!�҉�$=���_��[�8��C�26�@�_����`P2�a�m�z��*�'���:���5: ��фK��/��B{/����4[�G��� ����@�`/�'��^���o�h�L�p�Y���y���!zJ.��;�2�V������ׅk�J�Q�L[��x��#�Zo���q_���^��dyyy0;w7��7AË>Ӟ7��F�(h����~Ե���4SnӖj��<Q}Nϑt�$�j����1�?m!$̇�N���XR�^z]���������m�~�����V�Ɖ|`I���2���\�Q��Ȇin����K��x�\Gqx���&�眙�\�S�#�^�ݽ	�v5�/"��������#�s��O��d��f���KF�kAV�����5�����fp��a��A�G�ɬ��������~��m ��US��E�bY�:4�Ėj��c��ש�[�\D�%��l�l��tB.�Vl�6��+�����« Oq3e_=K�YD�7���ǫ�?5-6�NT�.4�7|���I?U㨮� }S
� _F͐�b�G�'�~�1\��g����`,��__�@�����}��Z1��E-��95�Vz�#P��v�	�XJ"z`�3dy;���E�*_+l;���*4H��i^�d*�ڵ��@c��x��L��~�/�-��Y��U ���ce涕M}PY�i�8��fU��'��e���V|��3R����]m1~�i8�#Y@�F-�o`�T�3(OYi����@��s�B����%\�k�&��L0���a`�z�7(n��Y4����T	�	]!��d���z��WR��5�����ޛNXr��ғ��	��!���.��n87;<Y�
H�x�%w|��)��d2��c��B���<S��C��&���̉I(����ګp���?N!���2�?.�/��%��j�&�"��e���{��a�d)8,̇^�˨Gq��V*�zQq�h���Զ�|�������l4���gQ��p��qͳ��ݯ���r4.����U�>�]��>���4>N$�;"y/p�Csi��n�L�Sh�(FFf �J9EG�r�Δ�H^��=S��"�`)�y%�0e:�'�LU.��`ns���.��켼����E���\�j�A����Q�diI~
��<�c8Q�4n�d�4gd�m�����~ݟ�g�;�V����S�����1"�7�E���i:XdX�$|gR1�Ҥ�͆1�X�4*�P�6YW��az	7@=L��f�۰3RW�/��Z7ĨF�w���ݻ�����e�B(� F����eUǽv?:��m���]wCy�Gؽ���1��t0����c������˖}���(ĉ"�X�#e�S�E��"9/
�&�$�을�MfֱGB�������~���u=��q�k<1�rWh0zr=�e���y(�
UE�|E �EvI�߯n"�͚�ZJ�*B$g�����4����$? IP �0�B��i� Q���>u����Ϩ6-�te���Ak�&U���J(CE��r�/(�J��ZJIW~d���
ZHk�6�!���lo�sԊIY����J7x^H^�cGǻ���:�̨�/?�R#[�yyy���#"αz���H�j0�3�����4�tL<�C\��̈́@pFY<vrR62�p�X����C�d��y���^ʐ������F�`�ڮ���wA��N�ֽ�$�p������v[�uʫcF�TTH|���|����)"�2�G��"�lM889�ش�i�7G3�ʳCz�l�������J���v|W�ԝ�pO��3�`�� �Z�T�N;���2����ϡFFF�6 ����Ծ-�ws��1P�%�-ӫ��ǽ��ÈJ�g���I�c�6�	&�r��/qz�͹mA1,kuww?v���+���Z)=��kq'O��78ˤ^��Uj4���KqNa���B��QFq��)���H�bB�+�8~r���h=!a�U�^���&������)Rk,�����՝!w��PU���B�ZL k
&;2�^��甔����Q��q�8�y}�z�J����L�B�B�l�$�g������?� ����>&���aB��y�<�;��,L�?tD�E.7��a�@-��l����(�/����tH�d��BA���ջ`o��S�2~�#��Q��ޏ?8�����#ª	V�\���`��Oq��*�n���r0��8�ϴ�bqJ��퉀;��`z�_�k#.l��v��pT��,�l�i:B<����(�5Z���k�urr��m�mL�����.�60^���<�����xw�"S�'qpW���ۡ5P���~XI���̷���؀,	:=�g��0��g��no�� W�:??��?Ĩ���������[�eo�ܷ��G��lgz���gm\0��	*%���Y�/�Q�!˶eh����ߌ�Rݞ�(m�B�e�:U�Q�g����(n��!�t��j��ᢦYZM��
�?�1m���u����u၅�9�#�j�C2��0�9��s�
>(��ɶ�?����,Ė�*��+e�^DuZ*Jr����-.��r�7��jZ�4\IZ_Yy�>QI�/��?[��AѬ%��Y#w�7��������t�>��]�SXx����܀5��)�ě�����<��
V��3}	9��o%�#p�Z(֔��gF�pFO>�y��r���1Ek_��~1���D9kF��R6U�d��_8�_>�O�OA��WJ�6A�1�wT';&-Ji�^����;��ml�������!;;;���]����vhvD�����"���l�M<�Փ� �˫W�γ��lN��G���%]3���.���6pS��ݛ)y�@��Gv�׀N��D]C��)ep�ƨ7��+k�5
rr�1w1�Yx��Łw%��D���?��j*���~��P�o�8*�)2)�|e����H�H���D�O�;`vq2/[N��d<e6y?�,S��T��Yj|�w�\��W޽B�Q�{2��볰�}�_�8���DT?������Kgx-�珋|ƁZ8��ElZ���/!�M!<�L|0�"�	�W���)-�XU|D���sqs����+x"�O��HOa�� �ۏ*�����[h�L9H�m9�v8ڪ;J�؟N4�66}q��~���V�!t��p"	=,q��Ue�/�|��Ͱ��)����C���@򴔯�d	��r�H�� �P|&�K��4Q��l╲V����Ӵojj����p	S\$U�J�������tۢ���L��H4y�d����-�Z����V�:��h�Iv�\�I"s�?���|Q����#�x͑��%ʐ�i�kkk)79�+�&��tt�u�NC*����ek��o�H���N�l��� �����n������H~J�.. �t=��,���UJX�d���c��E9�k����4�	`ԤUl�nB$����5d�NN9�چ��"�jcG�^�|R��<v�c�}����eej�H�8���:m>h2�� 7HaL�	��(��~����䗃?�r\��5��(���AbMq-��7�����y��'4���Ӱ��Mۍ�z��ͮN4g�r�A�%A��i�Uŵdb�-N�Pk����hm/S���5�Loc0zZ}Bu�pZ�T�����Fl�d�?U��Ou�O(�d����d�j�N����x(��%�|�|/����%3SGD�,��rԬ��E��!����*@y��̭���y)&��v| f�3�w�a����������b-�A�	5N��?_bzy���0=:zF���aMF���x����)�9��	��)>2�
W�����3�R�(!�:�فؤ.~tg�sߒ��F0[T{�i��	]S(�E��ܖc̪I�LR��������񡎭��[^�e5`,+[�pp���)e�xmHi�3Ŗ�8�
�����$���#��H=J��$��[��l�$��,Fr���3rӾ�J��vmޓe�M��gas�L+�
��`�}��՛��n1���.S�n�����GSy�a���m>�~���Vr�&L�̛C6r�/!���_ �ԋ@�bC�6�M���
Lξ/楟�,��.���x-j��ŵ�.���`�9�51�����t�8~����A�P\[[K�����d���%�}g�ڟ	?�B���m�ߤ���}SEg�99�|�𘲆�c�-t
���Y��Oי�(����ՓKV(����0G���Q6E'���<!���Cw���ғ�=p%~Wz.�p��qvۂ.x_Op�T��u�b���U�9D�7�PZ�t�.Q��a:D2}�Չ��bff6��¨[h�j�����!!�33
5�\�mz%��4��� ��=�u։�V����{a��Ab�z�!{��[X疹�YP�U��&��/u���R#��%����È�����f(�|0_S쇵d~�}k������:�!<�P��ZX�/wm?\?j�%���XmN�}�j�G�S����PgN��V�P�_�8=�%p��$s�;�������<u-�G�����̶`������T'�U
�j�6�������U�?�u���d4��I��:�'�4f��/��q��m�ǲ�Ĥ�]��1�M&��殃.�Y��l4ä�b����[ܫ8&}������U���'�b�]�J
m.��Ի͓���ɫw:=9��gF���S�HK�KS`�����"H��w���iA$�[��>IT��{z.n�xDd��L�ZP��o�U���ː~�mIfۭ�c�,�K�v�Q��W�M?l��1�Be����b���ﳺ�^�����R|4�	��y�]�?�0��{�u�x�����~������[N"{��FD���w,c��������.F����9P'C�9��4N��9�D_�}c�		��oL®O��T�As�ql�h�)0��+ �hK9''�bM���ڤ۬pp�9���7o�SjݙHCK�Q�`��@:��0k���I�O�M�s�����Q��?Uj�:�¯��^zaL�����Ӂ(���I�`���ϰ	dihMH��`D8�JI/jl�~��RԙҠ
�˛� ��71c�{kB6�@�$Յs��Ҡ���ݺ���,��F���Y�(�nOTp_#��?;1F-���&���'�w��u�-H�
9[Ѻw�y�z�?�nF�a��ni{�O7^�?>>�-^�'*�J���#��2d�aK̜(l�QlR{Bw�;,�����@r�2E�|��N\�}>T�.�5N&���j����oK�֐��_�XrW#~U��Y�U1���^ H��|."�}��naPXZ��Sa��F�A��G�D�+�T�Lk�������K�|=-~���e�]�w�`"�k�;9�j�
��b˒󮗳k��0���O.��v�_`��r����J��FĽj�I�1��!jߺԗT�c@�Έ-�9{D��K�*������U�d:=' !�Z$��_!�ںv�_i�F �ZH�Ӽ��M�Az�p�k�C�*3�J�x�}�9u�F��=��v390����7�(���Ą�ɒ��\ �E�υ�{$�\Ar����
��*7lͼ��{��$ZZa#��vV�ߴA1���ѷ�p�"u��"�T� �e��.��#Y��=7ND#R�¬��gύz4������:#�.�k¤�.g�h���LMu���ܹSk2:E<���_JW)f��M��~�y�1O�w�\|_�!��H)JxL��3g�0��������3��9N<����5����"��%��58�)@�Ӕ��J\?9�j�=y���<n��r�G���pHaN�ǁLq�2Ѻ��V�

.�O����\��ygi|��wM��Q@�L:��*D���N{Ad���E2z	���;\��)����Q�{9���$#u��q��\٢/*2ԕ��X%|�v����9Q���-"��i�`«�d&ҦB�����s\
X���P��s\��!&���Y��^�(��I[S�w%X��Y��u��Rլ�a=LA�_���*X�R�Z����Uf*Y���ߤ���p�i�t?����ǵS*�IS�0��զ�����~�>nf{ v+(��?��ؗ��zI8���^�n�#�A�h�?E+p�*��ZO�zcC��^D�Zj�[��Z<���B��
_lT�49�sQ~�(���Q�O��)C�(��}r�Y�M��+�7.#��bl�"���U,D;��t-'�ȏ*��߳ �,<�z{���&���_Ǘf��Ėo�4�{/*�Y-�\�5�nY�F��ތգ���=�-��J�ۊay���V�������ls�����k��X�[#q���r�_�/����Ц�@D6�d�cZܳ�0�/�Hp�67KRU���+i���a�#���-�bא
�Bf��Ka�>��������&ƃ~���p�vX	��7o���!�G'�1�d�ϝu�i�ɶ���Y$��)��LG���t������u�/��=c�>���<�����_ZV�Ü��f�΅�]a+i͘�Τ�-Y�D7�cu���.Z**��d��'ф�ޕ���O��	*�+ZT ��b#���M"7������ц�[�^<�����\|�ݷ'��'�_�~��/[�X��Pܦ?�?!'��@������8e��1/Z{��q&nN M#�\1�������)h���t�����WH�;��D��#�;w��{^aZ����b�!�B0;��2p}�����4�>�s@j���a�84[d,|��X��ߝ/�@�z��8s{K\�	e���7�L��ޢ��2�����X�'oQI��ӻu��Kb����\R� �[?ܹ�P�>����"�#h�2�i�����#�w�eI���#�!�(3㫦��]������ޡg�3�������������.�}���p�|��=�n/\=
�	:��.��?��>�y�D�}����v`����?�����_w���ՕMp��!Z��B��]�J�
��:z(T٫vs�㡺��?�&��-�y����VĚ!�o�~���)C	�&�a��
��«��j�?�]�j�{W���	'J�8��RI��7�6��7����%�d�q��崛d�����4��3�:��LLLf��W�?ʫ�ARA�̊s/Ėw������'9l�n��-��S��>�J(�l�c�O����Ӊk�Q6�0��@�$��}J������3G �$/w���I�Svh�a�Q��gɚ՚� ,,74�p6����4��W�ջ��;��I���&�4�ٷ+++�����k#t�H�|@�]��E��-���S�:��#KA��׎ݰ�t�W,5!Ĺ��%�!s���;v�K:�D��ͯ&�� �;�n?S�!�
��Dũ6*�p���p�CFN�Y4��6$)���)����KZ+��f�ͥ���3fKG���:���G��MO����7�'q�:~���N��1���bC(��<H'�ԗ=���B����qmueRuJT�"�;�`x<�7[��~�fr����	����9�+�� �������ی�Q�p��,X]˦bRF-���g]s;�v��V��g�1��"��!��bU�֖p
<7
�Y���u�<�*���M2{�������� X��(���c2,K�ח��1�Ml���� ���Z����O���,���TD�?���$n`B�5 d�O��]��~e��uM����X�&��6�%/�0H�6J��6��G���x����@�`i�^� �� 1VWG�v}�|�����jv������~e�|�����4��)E�h�*֫p0��q��xq�:��]�$O$��~d�.6�-�����
!#�0�Ur7�|�L�Y�F�2��抅p�L��88^S�������gԚ"��lL����c�!���5m�iS�9&�[�ߪ�����N�����E�.Yn����*]�= _x܀���cJ���dbX������`� a�ȋ؛>��Z1m�������B��h:��{$�PM��"15��}�.d��捷�pRm3�����e��#ٶd��G\��:�m��@SO�?��".6�{)`���@�1Z�^jI&�z>���C�YE���@������� r
��B���1��B����FG�P��7FOF��5��kuꝹ��yl��7� G؃����ሃ?�kjf,�����jrЂ��f�C�u\TN. ����\��'��p��12rh����_�~�c��1BX����Fa:���k�_.�\�b�+����Ǎ�HQ���:��g�'p�pU��&����c�;	�D�f�њ���qfv�ʨ��kxY�o!�����ҙ��LK�7$hg���ĈW;�Sg�ed4�jaG�F�;��v�+���C$߰e&��-y^p�um�1=�~:�22Kحw�Ո��9����K>Ӌ�[}�����'�ڀ�Hj�2�wfj'�ff3��LհQ�K�~"�Fv�b�Icw	�_B�՜��n!~&/+{BM�[�v��ۣpd�v=
G�~��46,�|0���f��?���%ڂ&��J1;AB�Jo�G��^�����q=A%�B�=�k�v�&��z��#���k����8��b�ܐ�6rU��^�	���o���� S�����r���}]|�^[�Ő�eQ�}1���t��QM�.��]��5�6|�@�$���Bjpg�@f۲[$����|�O'*�}}�FC�V�9���	����� ZHWR�_j�\� ��zռ#E  6�b� .0Xf���n�����pO�L8vo_�"�Wn�BUx��[��T���\Ծ�W��*I+ã����H���w}����k}��	��G���n_Ȍ(V�)�O����c&ɹ�ܰu������́p�3\m%��1[��Y)j�j�J�蒯ݟ����!�p��O�4g�Z����P���iBf�o���ņ��..k�in
�_��׋ �k�H�	v�\��4�7v�9����|�V�D�	!{;��s3����4W�n i3���kg�$ߟx���J�	�a��?�H�q.$���}���9��t�x�|r���2ȑ���\*E���'W��������O���:�v)�bcc3(�M��0>#�G�����;|J�ׅΆ��zk,���Y@ՙx�ދ�5P�_A�����֩��X�l1�y�*W3&o끫E)-lh��O�`�V%�X-))�-���}�����ր�<w�isqO��d���	Lv��L����w^�O���Z�ekM���$U<s�M!N@;�r���)�w�B;w/,,�߃	[��;«�ڠ�=KPM��@�����������?���eDm��Zͦ����a�)S�����.�WD{,E� ��b���8g%�"Es2�A�G'��cl>�tB�:V�kmRE-WŇ��i.FV���k_�Ā�"����5RE�r�UOF�i3Ž^�9��4� g�_�7�N�|E�?z�(�{�J!`�T4XX?���\��OG��/�P���j��.ɯ!^P[A�I��#����,K�8@�6hՁ�
%�.��B����W5���we������Z�q�����j6������3G��׉�+�6R�s���`��a�;�M�|*�,D��">?Ċt,��Y��^�2s���?�a0Np��|�a��L�����q�i8�$�)1TP��щ ��;ї^u�)b���#�@|-�,m�����RM��?%@'� Y� ���=i�����,���q�w_�*{0���"`f�U�e�?A���}łᚚ{I\5�[��?Pxy�� c�ɠ;k���@�d���}���n*��~�JfkZZ�G*�>/�`�����P��@+>Bӈ���I09`G���q���I����6O� �x ��;����{�c0K�������a�J�(���X���(���
��I��&v��ۏ�B�[����>�K�RL�j�^W��L���|^Q���Z�r����^�a/��qw��@�[r�8�1��'z1j|eu�Շ���(���ӫH���S�A���Q�F��8�
�ޒku���;ARE���B-�0ynMs��v����#��Ha&8��Ӹ�@0;LA�
]�Y���EWn������I׌�屋ۘ![/�X���B�H���H�IѧdΉ ��������U�A ���%|�S���+�FFF�DU�r�����k<
0�v7��3����5J8c�b	h4b������"�O�� ;s�G�=��}��џ�wS����x��c��$��;�a3�y�%c���"N��=���A���MΟ�����~���}�x���Ɠ����"2��put3д�\\��h͜]Y'Y�jh��_&�N�i��VN���m��8�/I��|c1	Զ��!��Ǌ(�l;$�:��[��x5~�{&WI��"B�p��q���`IL�����d��w��6����?ɯ�ЋE�G�ژ�<:s�C�4c�g6�r�՝&�Fg�~  +0�h��@�I6��C���6,TaD���o�C4�������Y#\˪f
V;�Xˎ�+n|��N���@.S.�fĆQ�e�涺sD~��M^̻�U;(��0��S?���h���HZ3�$s��N�F���'`K}�.���b�^�h��� �$!)9��' I����K�h})A%+'�$����v���l߯/mT|ЀoF�����;'Ē�.B"R��ERj6�-��G�AaR����<��z�j���S��~��Çi�!6ӗ������	:��[��o� ��ZZ$I��Q�7j�66 h�">fKpY_�|kf�ퟍ7v��˹����_^�g��M����뒥T� �����$o��ݓDk��Ti�ϏK]�$��1�˗�\L�јTZ��'vvh�I��e���Yo���5皸Gx4��i�*i�F4�z, �"KJ�
��{!3���td6�$��7���C[��R���J��l�7
A�o߾����˔V%�\s��՝ �������u�+���K]�CE �i�H�̭ts��mf�5#�L[%X�.����:�t��Ep�����^XS"���7Lא�I*��R/I߶Rm����9^�s�n�Y�kΟg��Wp��,r�(�^�Ҍq�	�G��(��3�1������گ�p��cV�}�FK��X|��J��#S`OKO��o����D�/���������1W̟�[Yw��b�� ��$�+�o���.m�S-�QZ�X�*yq��C��F�V��c\/׮]s"s�x�\�\q;TG��Ñ��	�Pc���/��%D�M�--r����n!\�7���D�)"�80�ӷ))�}� R������Ĭ������8�R��xu��@*p���0��1ߙ��i%d�ΰB�"15:aI���~&��7� װ{/�={v�%�A��ݬ��n���oz�k���q�Y6ac(A7��=�<���3���?C5k3h��S�4|� ��D�IvN�fY��ЂW�yY"[�I��;���C�?^�U֛:C�	��"�k�+�ݖ�����ǧ�O��I~Q�8���|Ѐ N���re ׉¹�T|���T��A�]�����{q��s��׺�]�˄5{L%uɻ�p�>���3}a�#�2�l{�f�-I��>8����-\���O�V>��6��\Vwr���u�%�1��7�1{����(^k��5{�v3��Q�З�ͧz���z�6+�P�Z�$������׋׊����tI'4�^��yh.��0�C�����2��0QM\�OQSS�5�� 4�C�=gHz%G�l�d�R�]l�׳���}˒?��#?�k	�vߗ��p���eE�]�ʄ�Ʒ���os���|xVF�0rN��5���N�]V&fe0"ը�LO�����L<F3K����S���d�K���1��̣���M���w1��o{�0H���+;;.�f�]�r	>I�[���JF���B�C<�����}��.�i�w�777��
���Qf�6���M�N���/�Ӧ��<�{��;m���	=jزZ�'x�t煿x��I����S��7t����7��!����덆�{�G[����0J�����o䐗t�VwAe�,�?׃�9�/�K�fTq9Ae��<w5�}��&,�� �~����rY�w��BS��j� �����O�@��4	�xP�ŋc��Q�]�b���:�L����]¿�����KP�K妻��ԥW��l<Hj`7����ի�?�@���~��[g�i�(#=�d�a5�^�cŸ�Ѽt��S��b!(�2�3�G_���(ġں�:\�ɧ?Ǹ����+�ᘟ�q�A<�***�:K���vhF�����u�F���������������ѷt�ݵlmmS�$I��nT;{�������
`����Fc�Zq-B)�k��2j+|us��\H&�X���x��xa�O\��y��Yݭ�=�#�����2]����O�DN2�,�;+i�)@���p�� [�f�����,��P�8���Dw(��;m�����O���>/�P�r7_�W�:%���c�I�S�&GG�o!d��EECxf�|�Gu��)v3�d�b}n>�1.|�t�����Ƚ�������*K~�f� �4@��K:�!�/�{��C8��������K�W� �՟,�od�O�Z��8<���gY@*T����u̝N�x|���V��F��kYN�H�T1ź��@�6� 
V�0�(�h����d��rm����&���}��/_¨Kl{����BKp*9����U�q��|�O?7��\_wW'd.�r���v���?�䧷w�����ij	�Io����J�>���!�tqz+�۠o���%�?o�L}��� s��+�{Ï)J��N��
:���r��wxLŒTM��@�Y�^��@��cm��`�ER�"�_��2^.����$���.�!d�~j/
L�e��=��kW��������}~�7t�s5�~D���t��c�E�r���'��:�w�Oܼ�G�4���wf�ww�L���JI����Ju�K�$�}dBJ����.���_�)U`q)�����e�����Č�`��d�ە*���O�z����� �^zܨ`��ѕ"Io�pk�=�~I�}��΢�2h�����T��G�T�����V��=D��f�C�%�Ηz���	�����Ǖ�����������ٛӘ9�X��yS5���f_�:U����N)9�a���ӽ�;��W��^�6/?xAL�װ�����q��X����¨�~�ƶV{��N��E�Aj��D�)����T�����H���X��at��y�:�)V�Ձ�䙰�\>�ۻ;sd����D��Nn��՝�N켔1�,�:�I��2\����9%�I�����~��-J�ÓC�Z߁x�8�w8)��e��%��.?���ʜh}��B�,���GG�'O��:�s���xC�_�yNV/�\&u�n�����x�<�n��aK��{X'��l|��Df���.ZF�W"-tN����uv��Lz`Xv�N̂��M}��h�ikx�U;(6�M��^(C5�0��2P �}M8�U�@���� ���vȨН[��z*�����ԓ>Jd#������I�����ё}���ѻ�W��yg���ǫM����������T���6䈦h�m���~V�9�DD����.��\�Mu2x:�-[)�o�۝��~��W�斖�bI�,���,��`��$�£3Y��^�-"����R�￮s �d�
���	�ڜ��I���?�p�o�k\��U�~��=0^�8|4�\ �Y`0�M!�>>��0�,I ����_a�~)S5ʍ=�Z�9����������+[�yu���(0ڶf9�U�Jݱ��8�����Q�4���Z�^��A�g���z;a�� e7$�'v���?0��#�"�=~���(���)�a�[ ��'8x��F�a��i�V�6&�m��@*A�=}혯���+�n1N�	�iY�ϩ��-�3Vp1vq��^�^*M#��)�rW��%�Dp�zx�ߤn�����Q��_���	b��E��A�{ؙz�E���'w��<�$&*Z.�3�����������|�+�aL8���t�z�sps����QjlJV��8P��Y7p��m����b�����B�K����:��Z=�k:94��_W\������T�M:,��ro�����p� ���uX{<�T"E"��	�5
3�#��PA'� �bk�w���WtD�(s����/������fN���"�߻r�g<3:*i�VΙG�{8���M���+�K��^������Ѷ��/:�#"����YfbV��x�f65���G#��ʦ�
z����/�fi|��\�6��i���o�U�~FFF�-�$��&���V�TQ�-�/����M7ϛ-gLs���������8���q�
q�IO��ޭll�=^˹h���i���C�s5�	t�硨��y�i0e�l|�$gH����E�~ٿ�[�{t�*rsR���:�����c6�Q�Q�����s�<iKH��%����A�,��@�|I�`��ѷ��uq��:��+�z���+�ϲrT����W��
V��G7n�q�,�����z ��E�Y`��s��'�͈߰Y��9�����������t�"����	
ee�-Af*�<7��4�ϓ�H���қ��ri;-��Ӏ�J̛��Yg����I�3�����&�v�1�nڐdl�T&��%R������,�sOW:���?�#��<�%�6w�C#��^ؕtk��Q$�����((�ܓ\�xF ��y�l
����1"NҢ��z��eR�MG�d��� 6�����gg�U):� ʉ�K �/A���l�s"��^�#k1l����~��0��;��9��w��w��4�W$D�������#����gLj�����{�3)�^	��[~ܑ��4H�l!?漅��u�'�Cr��Eװ��&�f��������I�'�T���;_���֧�cN�vS�r�����Օ�R�߽e�k\[__��}4U��)�"ǟ�(���W��i�Tr#���u/_��~�����oY����#f���������n1�I�U[L�́�,5I.���0d�I�Q�^���.=Z���*u,�,h@|��	G4)�ē���igxG��J���M��<�l�	�b���>�ԓ;�~5Ů0��8z<@5(]����;j�tw���W�D��6�c������{��:߮���E8��<�]o/C�-�馸xs����UFjt�s��T�(z�K����W�|��/R2��r-��A�R���R��W�t����_�t�6����@�'����B9> �ͻ�9c����93�ٵ�b9�?/T:�vV7��z ]5���'$��Qk+0B-?���?�$��)��F�Ӧ�� ����Ue%T��~	~ED\���^��x�1������(a'��I�t��,k�0�/�Q��/���~kOvK����aW����r�V��}=^=`�(P}16�,�ְ���Y���h����)�F�t��)C��Y��C�H(�g��i�2b-������|��}ʔ����zՁ�L�3ͬ'�>>�~ݺ�g��EG��ޞ!Ir�@ja*��o��2g�$%%[J��g7��:^ל����L&¯�^k�188uok��I�fM<//���ץ]���d�M!�co�	e�����m 9M)���9��8����5��(�0�u�:��(㎙G�7F���2'U$��k��#��c��G�el6e�Q����ӵ^[�<��m]|N�/��n����#}��ȃT�ɉt�
��^��LwBc♩�2�tU/�q�I�4
�id��#��u�j����qB��F�ޒ����oRD����Y!�kw���m=�~���J�.�x��"�v˸���ݽ����~�D7<�l�[�O+E'�]��/���;���I��fs{�k=7
�j��[��3�Z�zs�hWm�w:��	nw��Yݟ�QU�tK���Ѽ��W�%i-���l��M<���6
2�F�8�d����
��G�a�/�&!�%U*/]$*���-�\���`�"���2�W�M!u��m,	�R�q�rrr¹8ie0��E�u*����ƨ�皯!�<H���[��-�u�'#�lm���J������_�!�Vz��è��Jf8y���D⁝k�u���Lj��Ո���Yۦ����#���gI�*Ƣ�RRR�G'��vk~��e�]3(]�_����QO[��"�J���ei�$���9���(��|�aou���qce�ڼ���C��9�YS(���w�<�(/ccS|}�	���vh�ɛ��n����H�=r�����l��t�oD��,����S�(4v�B�p+�v\��%�6޽������������Q<���N�ɟ7k5"78�MS=F���爨��*И�<���=��.��,�v�J��#��L̮��%�o�|��Ӻ�r�v�J"�e�&���MS��� ����:�6U1H���s|������>��^)�E���}��w�rgD�t^�����}�/5+�j��f�����#�V�S`�!��ߵ�����%�w너�^D�/b��'<��I�����0	�ی~h(�����@�U{$�-��d�d�Gy~�A�R�S�	#k���ã��ϔL΅@`��!M�����ǩ��29�ְ#�B���=���Yb��
׷�ھ}�y�ۦw70A%הnVjݶ���O�+��0���5r"R�WT�����Ӵ7����ls���[w&��� �H��I������}V艒A�hp�^A��yi��Q���
�N�	R������ыQH}p�wW��&�� �Hl�\Rg@c�_MMM"�C�WW��i�g���_�$2���������D��?�� RT�{�pNnڀ�BmΟ��d�z�*ϊ��㞲r��%˧a+s�dU�_"�D���?�?�Q�%��y������U�M�����m�Պ�u�Zq��|�{�GYl�3b��,b~_�Jg��gx�Io�x��nWkYJ��헸I�_�e^[�z�'M�N�=k>I�jO�&�Õ���(�#�>�R	P��d*f3vʬ-����~�e�\D��x5SG�i�A�=.�Z���O��NNo::�ʻ��[���#M�d���'�E~�KmoȈ G� -��Y�����1���{W_���U���0�M��{��ƥ�I��|m�C�dT.69�lðu��?����݋
��p>���dŠ�W��lJ��0�&�7#���~�ۻ=���U]��x�
2zD�2&Z�1q��wN"�X�3�������<P;��r9�
��;P�ј���Z����W7�!��Wm;�kl)Z	&�ui�)S����}��]vO�u\?oZWp�f��@Ĳ~��t�M׮�d�>��pzb#�"�X�!����e['ފ��'���xl��g6� C�U틮>�s9aD� l����Ų%�Gv�~m4b�G��o�w���ʈz����F��M2>S��˦A�U�;t[C��ɟ� 
>���N����N@AHϖ�Q�3f�ƽ�se%������U�O�RN5��/ǃ?v���x�+k�6���q���[��u�\Ru�������x2e�����e���4�Q�;�cG`�ｶ��[�3��_U���ʣ�Ǆ����yAܞ�

ݒZ����`�����sw�Y��;Ґ�ܤ��ʭ��*���!���^"�')�>_N�X�tw{��P�&o�ز�|���Q�__���}`�W�@�e^u,�B�OIH��,�/\P,��㼃[Y�tj<�Fc��h�H࢈l�6�J�<^3S��m�����(=��M�p{�/�ؿ[�sC>E��A-'H����w�+��/���2}W9�X��b2��e�O(��7ioдT�VVVn��$,d����$Y�h����V�4zA�%�&�3���վ�f�]�p5R�I#Ѻ���M�Z���l��ȗ�®��ݐZN��<Y1�W&fj�.g}��œ��2�w�WmL�ϛ��[p�������S��I�*���èL0��s}��k$#nYc���-�����^�T�2�4uU���OV���V�Kv��%�/�D�s��q���QM�<��z_����_,,�Di���D�࢟���].ƾ�V绷�)��C���RU��!L0kD�!,ȿY�7�r�����1�\CO�79�5��}�o�>V��f������:�����jLr�5f*G��.ޮ�R�d�泌'NLW��L�W�V�!glPP�`)����{�ö 3��	���]���a�m/��d��? ,��J߼����Qa�y9���f�7������W���L���Ǐ_|�"v���P��M����#&������$h�ꦮ�����>��ϸĺMI�n|�����@��q���hF�=����9m��C�t�~�w{����K��?��<����"�lS�2
!�B��k���c��Cv�4(�d�&��}�R�d�!&K	�P��	�3����{<��G�s�뼞�9�ޡ���������;r������8�RU�t^�Bm0�/(�=J�����������=%lR#��l�v����p>uK>�0�?>�=1J����ԍQ˝!�Z�Qm[샦e���P�*��;�>r�lH=S��q����W����?1�}�;�Yi\9�3c)L�<�:367'�קt9S�[pKe�&�#��|��?�����9��b3o��l1�vz,��*��$��T Y����0�Ƚ�b�Ll�����玲%�[�ؼ��mC�r�۪��bBO��rڮ��:.�H5)�On�3���Q����Peh��uQ�H�;�S&%�����~��:c������^'n�to��@����SM�݁"�̜����B1\ˆ���6�s�`Z���� ����L��I�˱�[M���S�큢��#ر"�[6�W�Ӎ�?��nȱ.���t�٠P�v�l�.Ec+]�Foo֗6G����
g�ȳl|Ue�
AO��I�EjY�g���ӒL��r~1"U�X�� OF1.}���s
�f�������[8BƇy���F?��'��/���u>�"����e	t��g<Sm>!^yNJ���N�]7���f���k�M��NC �e�A��{6���uڋw~�;�s;v��ƃ�/Ay��S��F����/=n��u	��kf��kP�XiT�Qhv��˗eN��drI� ��L/qtF�.@>0�8������6y(��ź?qJ��mR�V�+�����n�,�����":�p31ޭx�T+}W��RFR [�$�S���#��8܊�4�#&��ht/��i`�h\��_��~��Q�>��'#�WWW�Vo��>.��L�d�" ��A�T@�r���`-���llK�M+*E^����R���o�3r���NM850��0�Һ���6�
�O�%D9�3���}\��o��p�!�bhY1$'�RT���b]MP�\�%Ɠ�̞��w2�,v��
3����s�R�]~L�i�X��T�Q�{D�P�+抅)j� ��!:�Ď��tsP�{x�U��LT��_������:d��[��ɁH�Z�m�z5�r�<�cI�1B�I.K�Ж�iv���_8���J���-�Zz��\�e^�J��0�NU�{��D���ނs�튏���e�ar��e/*ڕ�|E׷܊E}[gy��V͍�����|1���b�@�;���5Dws�T�X�_�?i��D�����)��c���ܴyڿht�3b�C��<7�q��O�q��n)����s)z.����Q���΋~��%S\�k
;�)*��s;�>OV�p��VnT��L�Qm����+N���,ʱ��������K��8�#>�<b��ב�?kC�E?E�ήLԂ�'�����!�hx�;FD��/��!L]q	�Hi�4w�u�c��G�i�נ�4#,Ĺr|mw�j���Z��>�]]��|"���^8�̽��)��4u�\�˾��B0%��PY:: �$)	vQ�b����nc�Î͹����?7�{@��x���O�y�}98H�"�Jm�.�Az�����K�J�"�נ�}�h��0�K_�������v�z�~��]n�w�?\kU�Zb�f�c?"��73��X[ݬҌ��� v�A�#4j��b�T�^$�/��6ݙ�;��rN�_ܤ{��{E��F�?������$���,f�*Ge�Ĩj�I����/�Z��	��~�x��*>�]	�c��ϝ�~?��g�m��~�E�ay�&�s��+Zf�ڀv����#�i��x�$���&���e�y[��Q��)�sOZ���������$}�-�?67�D�������#:���X௽}||�_FN5b3ӫ�\��M�r���iL��="�m�9Vf&��*h���ܙ�'��K77��dϴ�,�~a��<��@���<4����_E��5@S�M���I7��Ď�k�E�����l���l/�4 *m�ƖXkP<��9--t>y��㍀#pK�T���>|`~��\R�4�|d^R���<�$~�3�����~E1����y�"��tB�*ٔ"u��:�vہ�N��;|�<����܁����c����[��cޘ�U��JW}1F�b�<c#0�3������2W���ں��p�N��ӿ8ط������o���Tj�Ґ\Kk~��X'ROYD�U�������e�:���e�M��������԰95��T��� f����������}Q[+
��������f��`���j�E���'e�[8/�҅��	K��c�����u�u��z�)-Z�~5��f�&u��7E��d��sK�5��Zs��b�z@׹ߔ鎵{}�W���O��IQ���2�ډz\3�8�x6����3pd���P=@�I��/�����2L7��E)6��?4��瀅�:9 �ܗU��.�z�Э	�e�V$-*�_2��<NP^;�vhs*/rp���_:�7��@��<�&�(�LÜ�\�{���A���PE�Vm��ƨT�B���/[� 8����I
d��D�v����I�^e��d��`l16��u66��`�Z.>�XIƅ���ᓸ�;V�nؓW���h�XA/i&�%�k�wg/0+KL<���-J���rI��q�>C ק2�+�-Q�����:����ERM�W9{�.�8d��:&���^:0���4���!u��w�� �W��e�����B��
a��.��"�~�ʜ٧&,���Xb�h���|N̋o-o7+��lg���^���F:����1�i8��x��(J�%��%��[�Ҟq�<�!��tn'ӫko���j���"'q��B�tJ�5oR�s��#r��W�.6�����:d��v���꣹y;�ֆ���=��{|�>��X+��~���E�0r������l��c��R��k�Om���\�^�sMS7D���%n������e�N�t��u�!���+�hw���k۔o�d{����'��֤�b7�^RΧ��[W������9��_�zU���MQ�r|Ϸ�|�w���Xq��J��X�_�f�,%��@�ŋ��G�xc~��qU�Fߩ@���܂&cT�̀f�B�Dgy1��_l������Uk�_ȡ���kcla��;���y��L���h�I������@�gb|�e]���LKrBO�h�tT�V����,@>�t�9W��9�����N�I�/�b��"x��Q�L�d��LĹ6@�$!��_�O.'3����j�K��K!`M���|�*}�ܐ�﹞�[o�`ݓ �|ti s�
D�s'�P;�����бq�hf� �j>��o�\%���8"�h����i�s�NI��\�_Kؙ�C�`��*�ߓ�鲒��;�x�+����*-u��^�~�����a��&�b��z�]ThiV��zE���
��"�eh	E�nĥ�n���qS��M�^�N����!�5���� ���&�����M���ڭ�x�֖��бq�?�S���cx���@+�
���<|jT���c��Kj4�pD6b��_.�g�q�{[j��H`n_QPկ���A$��c�y��H�d��˙%����*����f��(s��KN�h��|��b+�<�������3�5P.�Ɖ��׺� HI�.�����r੍�^�8]�� ��4��f��l���ʧ�Y%,d1��/�=v��9�����o�$�����w�����:+����ƯݖJ�{��.s#[�
��{�uA3���O������*��_"���|�{��4��|�K�����#��,�(������j�ҰD|�Դ���]<��7w����=�YY���wQE��m���nvP�;�[�U6���� ��.���Y76Ɨ��_C�WW�z<�}ѻX`V� �;��	 ){� �6Q���y�R�qaB�x�N�/h��Ў�8�5����5vP���77����+0��s�K�]�d��o9k���|�f��ϟ���h�Ɠ���y@x�J����ᐨ�ڄ�KO�^[��Y�߬D�;�vc��u�'��ZȎכ���lH�
����C4�%0>����s��~��p&`�(ʹ����^�\@�x�u!<�\Üh�F��j�[q�y����	[�a��{��)E��ģ>��.��e��@����T��+YEV1#���=�,��(
�@����j�~�Aa�p	!��+�=~�+a��
�ʕ�r oy{Wssоc���T-BP�����X�lY��3dc�×Xm�6���Y�����X�%�('�@����駒��Y��n���M�<ls�zS���Z�1�R%�9����F�����<�66�%f&�s;��}� ��b����J�	���'/Jf�j����m$KYi����_&��lw���d��׭�Ԁ[�}�j�R�ETf%�":6���ȟ�Z GŒ١�O�4�6�/JSdc�$Ȥ��]z�SW9��U6!�k�wO|�ٿ6�����UVBl�m,e�%�+y���P���UiDgag��j!Px�R�ƽ!�zR�WlRK�1�ɳ۴��=m���:^��G?nFh�#R%���������2v���7i�,,)�R N@{q����y,��*S������">�xnZznU+-�����0���y�[%�����\�&J�(u�rvNW�%�(d���r�v�ߜhj�X��&��q	�:���I��n����u��n��sL&�qm�3�z׽�������:�	�tR3K7��&G9J�X� �+������'�L@��_L�e��]DDꃫ�C���E[��U3ĒOA�W"*1>>������ �|���;9
��1�;E3�=�Q^]�]�z��00S���<����;_�&��@EX~y�>�u�Y^�㍋�ѿ%�I�΢�?�D����C���0GQ��.F�n`���w��_�;WZQ0"ʔQ��0�X1ɁGzչ*uC��)h*Evn<-vtS>���Q���f�K����I��!X�?�z��2΋�j�����ݟo���(3 ���E���j��~�ݨ�z�.ʥ�Π�V�܉c�r�܅�ݲ�4m��lRGmx)P�Ư���&���#��9+eY��VY}��i���<�҈����#��M�;<{T�ɕ�=�v)�?  ����({�9P�ۀ���1K2�����}�c6'��q��g�+-�9�%�1!���V�s�$�)��m[�>��Ψ䜩���U��� �md��	0�;g;2rIm.	O�3���z6�WPP$�K��.W+I�5����*U1 gH�X�O�!�
j�D���ϱ��9�bZ�Q��KX	��}�EN���+)}��g��I�_�Ĥ��CĜ)J�M�W!_�Rt�����h	�B��
�#�<v���j���W��?6���z��SsC�����Z[[�L%�#����M
r�e�bT���8���j&պ��7x�ӸyC@#���nB��d{NV�oJ}�ʹ�t�|����h������~k�Y�w �P�u�Q#�T���B����.�D�r�.�r������6�I揆���ٻʨ)3U�>�O��w��R���	<i�%}Ā*�#��!���`��Ɗ0!��F��ճ�X��Q%��Bd<'�����,vC���|dhH�� ��b�Y��ŕ��_Xթ�3H!e�i`d`WJ�z� �%S��V��g�qOC�Z��n<��bS��m-˺�>�{�0�Pu�oGd��˹6>?(�Dv�=<<<�����E���V��%FVќÚ�6>�7�)��\"E�Y>����"p����9�M%��#=��k�m���:=�B̕�ާyNQƅ�s�Ug	�tnʱ������~��~;�Fd��j����w��M����F������A�7C�/� ,�\/Ҷ����)����ڥ���fH�.	1(��^\��\�;��#�¢Wx����g�m��w���ڒ��	?�I�Ƴ@�O$M\�:D��Grw5����:b�}'!X��c��,5`\8�y�bΑWFo��vvv�w��&���C�僣x#3�|��/ϥ)v����?�^�����v�j523�Īch�8h��	��^^S���P�f���Q&�xT@��G�G��cm=�ܴʪapO������(&]�21��X����,����o�(R����;�K4�����Gמ����?�	�w�:�˒��^��C�)z�k��h�VPP��{���a����	�V��bm��x,�%K��]��E?℠]Ufہ_�UZ��MP��~�!P
���J��0õ�@"��.I���F��z[a�C3_W'ļ%gbH�A{����ϱ�5�s�;���q2�t�#�o���B� ��e2�GA��o��V��o�wJ��x�+�%�?E�R�Tv��������]��쭖h\�$]��*�4^R�wn�h�X��JI �����x�Gn�����||��a��,�%�7y��;�u{�O��k3����Rp,1��K��5;;��z�\Ǳ;Ψyq��1�e,��N�u�l,b��WN�� ����}O�<�pEƶ>���q�~����ҎR��*?R�܉&����-2va�A��E��ډU�_ξ�K|�Ef1 �D�V�CW0[�/���UK��F�cI�KG�'q2b��+ ���b����0�1۪���})�'��8��꾯����E�^�h"� &�b��g(��NS����6Č��;]������'�f�QJ ��?n��Z��'����P�B��']�t�7��)�%R��x��L��Z[��gK�c*��ﳠ�9�����W"��
o���(����5>��zG8ۨ����/AA�xz�wlM�U 5bǯ�Hqo�iC�dm݂�v����G9`o�}����Z(�G�dБn}��Y��:d�j��;�����.s�¬�l��8��.��y6	�g+Ɵ��,���XYY�)��f� i�j;=�/_nk�g�v�y��>d�[����/�5���"�G�Ĩl��H4���c�aa3�I����$q��>�Ȉ�ponLv!e�c~�N�k��.2�z��bg:^uUiP
��I@�M���"��<K� ,�,��6j�*�S��(y2��9�^A�S�DFF��M�8�7WV��v�C��c�_�@�� 5��5V/>T;|�#�X	^_�E�5b��𸏸cCA��q(� �W��qakM~��8L{3{�L��1b���V0?[�n���E{�oxg?W��O�k����F��+[���I#D,v���X��	St���ٺ���c]��W����l&�}/=M;��̾�O�"���WB��E��w��|S�_1�>�W��*-ċ��&��<\1��o�nƩz�;{\�h�S=�rs+J�AT*U�p����2��I/=Ӣ���o�])	��H���Yq'Va�Ѻ�Y�عSQ���m��O°���Y���q9���ֶ��ғ��;S��1:Wo,S����t��J��K�� �Q� }l~�K���i�sTo7�����%)p!�������}Nm7M��lK{�E��*��X�����N����W��2ˑ:����R�!
p�^'����h/�ѡ�xX�W���7;�vUƯq��,�6�H�g����Sb���;'~��y����`�@0O���i7�#+k��$5r�
x�6��;*�I��^	�C|��d���$@���e��+��"�~�}��xAI{��Pҿ�){>����ɓM��׵
�Sy���_���~m���@"�L����@v�c�t�V�as���j�K��;R��0��߯������%h�����֞�%U3��D1�16��K�ĭ�L?}t*9^�4�L��c��q���<t���R�ǭ2�Źl&qvL��Oa�ju�"����>��T�)Np�k�w��>��	o0l��ވs���Ȉ�Q�w���`���W�n���6}gɷ��e����*�8z��@�[�@��,�{<8�6p;�����0�J�9Ŏ�9H]���ߓ�́��"\i��x�_;�m#�V��$>�7��Yzwh���(�@�o����a�\'�mIRV�Gb��ڔ?jy��񊈈�F������8��m{�b4����L�i����z��,�����y�p�`dg�S����B��A�euǣ�9�߯"
��TAo>L��7˟Ά�Gt�`��܉�+�>���ֶ֚dw���ǯ���Qm�^��HX�Mޭ�z(]$B�`�M���ul��ݾYAڴ�o���֨���l�!�	}�a��Ӳ���H�Ӕ�je�'	kP�m_,��bT�e
.��Ѩ���2�#��+�)O�9���ךw��轋Qp��8вJ�b�L��0U�=4D.�;�k���G�`�W�᭮#��h�c�)�l]�5��MN���/��+P�Y��ʽӧ{�
B$����� �a�r&|���
	����Z8<��;��\�������q�~���V���v�����XeD�A��Y���j�ɑl�A�}P�`��I�,���o��[�ˣ�6���rm�y�*��9��)K��-6����UT8!q�1<yA)�+�GPpv5x��),5�J�p���k���k���K�'Ǚ� ����m�-ڲ+�]�˓$�m�+5�r4��w�d�����U���:Qa%���-�\����"2@n2p���	%����E57"�_
]��uZ��l���~)4o^G1���P��h�;��W��X�7+-@^ws��3˓|Ḡ*�~�T����9�p��kB��N�����dU��X��� ��g���=����A*�O���k� o�L�\���ڟK���DL}L���Qz}�"��)�<���S��h�>�D��Qg0��J^��\►��o��\��.5�y��|j���؀%5�T���_�;-��O�s�qط���;'��be�ַ��I�k�U�ڦs����D	t/gj����j�%;����G������e�q誕:�>��HM�����<�� Z�ԑ��4O�t?EǭP����eܿ'���9�T�|�)<}|��$N�B������n8�5��Q��T��m���x�Bvx
3��Y���p���C�8��|���Y[1��΁N~��pǛܹ�M��_�

ک�¹��[6���@�<�ԨV���GW��c�G��2M�_Еl *��߼rԇ��~`�ӂA/����H7P��r�H��O��v���!� �o2�՘o!�@=@z�2��9rK�P-S~� !��a�1��5>_-	��)sYEE�>���Ļ�=C�����-,�J73��&���rr��U�_S���_"����<�ˀk���+�-�����狩)Ǥ���G����_�|^�yZW�Im�� �3�?b�SP9j��&��皅l"�Ծ/Z2EϬ��E&,�v���	U��?ί�_�[��H3�+F&�es�ۃ�wg��!�-6�0ƺ�j�������u�WjDؤ�QT��ߧ�b�K�;k6_��,�9�C@�����l�A��0c"����V��-T������W��᫘�'�D0�s����
d?�\hv����7�R�����u²�BN^޳{| �t���J*��A��G|�9+\�M.^eu�C�Ӟ�m�>]PZ.c���^R=�h���r���s���;��|z@�Z�1�O\7��-iQ���}_hҷĥY�TQoQ�}�`��Uy����8��5S��W���|��^ݐ*�F9q�przFD����Y^�I���,g/*@��f�Rr?�_����c�8�	��eؓ��.k����q"�r0syH���A�:�s·��);;g�	�'0���u��,��o�}`V�Ay�>hOwEօ|/*����� 0�)����v��ZfkȤ|<`��!�=LN�Q�E>=a�Ὶ^A�G�������_9����X��$$I����eR��W����ω��ˏ׹m����@ ��X<���-7g9<#=|��5�*?�֨Z57��DEƄM�����Z��q��m�� �e�I�ѱ�<�ʱ�׏�;R\_/��N}C�o�E�
3|J�����������k��ny�`����
۟�=�8�g�?�a8-��+���꒞��
�d�j�9�����m!����waЎ�u�۽ճ�d)����F�r�Ҥz�Y���������P�����[�<����k��BzpN�'O��ьiك#�&����f���^0b�{��l����o�/�NĒ�'��!�eX�fW���lo鵁?��hEn�}_Cj2
����Y�PXM�5��W�8�<lD2ln�J%���H����6��oE��#Q\1g��wU���<,Y�csӸ��DTQ���NŨ5�W��y����!�p0�:��fq�0�h��|G���7����X�}�<�%��v�����/N��"�j?}��l�������F�];x�V�V�����{�뤦�ݥ��~�H~ߤ��WC:1r�� �򶰿�Kz���z}o�~ω�[�δ����u��G������Zlxsj�K_�7�����Ξ:/����"��gdt�5Ek�,[Oa��Q7��)=�S�R����V81|�'m[8(�����P�v�T�'M��+����8@��[;�\�Qر֧&(�S�Ծ��(�I��0��e���+��Q��z�����5g|����^_�[5�Z�3B�U�2?��_�:���v4�� ��!F�'����1Uy_W�y���{�Rv|@Kju"�g�0A�G�c9� ��?]����ʧ�.���ʌ�2h&���e��
�FnYTPU�y�ϱ��à~���S�FK�D��$(�Q�Aϛh|ZV��ܲ��Ǘ��\kݸ5*2�Pzݹ}|f\�o/��~�G��!�N^=�W�jw�TL�S����IA/���R�]��G�+b/wl�y���T�ڮ������o.��޼����HMT.�~�&�:f��6���Q[|LT�Bͷ����N�~X�t�	Yî�څ��S"uKE֕���� �q����Z2tq�/���34Q��	��v)�%�cҴ���e����|h�}~9N��-2^�&xr�Bkڮ��@���Ws�Y)WN�ƕ��h��d����(�8�{����N��׷�)�xleУ0b�m ���B,YO����󢏵������0S�v�5�����*;_��;�n�j�\B�/0j6�%�;�轒�_]������}���J@ȱ�::�*�4�t9�n���{��_6�z��_m��	K��ƥ�,���O���i��#�7E����#ɉ�o��V�%Y�����L����<KP�ofS��U�6Lj�ѱ�O��Ƞ�ѥ[��fil<����v���m?�<��O/���,�@����gb=(DP#67�s3-hL�����Z)�E�q��)F�Uj����C��)�mU��k����k��uC0�6�j�Y��:6%�A��vS�@(u9zUi�9:1�!�"���J@n;"<x�}R#�`})Եշ���e�����7@�h��a���֍)c���	�`*�J�CY��Ot���m���n����Z|��w��f�r�n,�A��R�ll�@���v��L�����L�B8c�p�����s;��d��)��޳*%�!4�H\6����܉cČ�ǁk-E���/�J��rd�%[�yA�55r��8a/�.���V�~e��k<-��2t7g��$���	��4P�l���$?N����^b��2E,$g�dUv̊��E:�uzGл��`kk�S<64�I4Y���ZIv� fD�1$xq%<�Us��0z��Vy�:�ɝ������gΜ	y8do�n��~q��<�USk<��')	��J7���\�KeSuܡH���^�����O�][���J>�y�2l��Aн�{����ļT���M���I;�u�twó;'�J�W,Ͳz�`� ���j�����}��:f���|D���[�l$�œä�����w͸�=�%i��S#_%J�nN�"�2v��w�KU�,��K���W�:���Z�Dv�+u676��]D���ru(�>=��'A�/�օ[�<�+
�����U�إ��L�������<�J�e�y)�E������*���k�pc��g�M�lMf�F��q.V���|yX������C/Ӈ'�K�x��<��v��&	��� ��^b+b�t�����$U�P6� w�N|xQ��>l�b|Ϸ�F,���	� �ÕO;��5S|<x�~7�R��_� R��/b�Ϗ:��Mߏ��/��j�{������Sh66�1)�����į&��
.�6ٖ���7K��|K>c��ģ~�r *�_h|�	H/�!�
_Wfڮ2(�p�U� u��ca^:�|�~�o�$zv߱�/Cw��I[{Ζ�%��0��A�vF�/W���_W������ �'�����~���RK�کO��Ύ;t�'q���ٹМ�a���utv�VR�S��ɼ�#}�!��s/ ����;�B��ڈ=<�Ճ���V�v(�7�pk�=D�ɳ���*7:����stν:<�+D(?�ԏ�읈=2�R�ʣgX�>�F�^)�#ǥ�kjj��ٷ�ԃP�+}\#�S�-<�H�V�C��K��U��E���%��{}[�{[��~О��x��˞�u� �f����;�WВR���%AJ,]C�_+gh�s����V�T=�6m�F+�$��nu��X��^��Zg��U$�$KPkUh���q��Oҽ�X�J�?�����.b���p������`\ƀ�jO<ʟ��R�p�����r�N��e��umm���.��Oe���i����ߩ�:����#�y�����k:��s�3�T�z�aV륮%%���dDd�7-^�m�U��Vw�/�gt[�~��C9������!�_m�H�S�tg�����Sg��l��ᔁ���
	�O��=���d%BUA!ƣ!Σ��I�%�K�f�%���9�����?�Z�c����o�z���"֨T�o��L�Z��z��brwh�H��X	7S�~��ėߕckoF�U��wZWF_�����)@��p��S;������&#������x��ô�@������s��2�'p
�"��eNn}��'�&1c��~&�&�q��/�J����&�*/�&hV�D��7��@�_8Z����U��3�Q"�������1g��"���K�Ne��w�D}栟�Vo�m��0����շdr	�J�=�qBBcؑL����\��{����O��`���L1��\yb~1���O�]@}�����8�+9�S'���1����H��$Fyq��c�,R$&q��*2~= v�/_I���Rsa0��-�w���B��ly���E�*�VN%3����\����?Q��	A�S���^�\Zɴ��_���:�Չ1j�#�aԠ�i���RJ�Z��8���@�
����_��G����c���&�����A��0/��������9Ͳ&]y���%}&(o� �
���1��@�@ޱֺ_�.��������yǳwyr�6�C@Q��DCBBn����d;��G]t�&��U6m����tδ��O�K���c��.��u����;��tP$p����g� (��CX�cĠ �*ωy����ㆻ���M�##b������_���z���d}��r��{g�����g�J��wϸ�/��s4��?uΨޫ�4��U֦d�ޛZ)����ͭ��x,��K!�H5��pU=� ��~�fI�(u��k�%t&��Ŏv��8��<�9��g��;�Q��r���r��[Uq������H$�\/(F��\v\֏��ʿ��N��-+��\�����넳���f����MO�*!AmΗ��q��{�ص֗�F��ͬ����95�.]��1L��5��k�����]J�rpYw����IR��e�Q�����.S����Н���I�)��������ސ#XW�%���m��:�Z��m�7+�R��<����3��ҋ�_/(�I���6�,J�p�ҖRT/]���VoV�ud��f���{*/��j��]{�D����s�!�w]���*	���,��:��y{�����nػ\�u��H1�H��لy��ZiU�nra:�»�G|�}�V�0(f���[e�a�=+h���	 ˉ����y�$�s�u�⟧��]��s[e���?�7 ���<���X?�Yp��X�i���5���+�2���볈�j_��7�a��H}�����@�=Ӯ�7��/�W� fj��>�����赧��{�MP^g�]c3�D�tl�F���s�� ���wb��s�M�ݸ�z�w��ۀ��\�N�~�X�R��$�mM!�]@��p�N ������WZ���jo�FQ{hkN\.�x�w�m�K�-0g'M%�������R{a�~V8������E���N ��l�B�ߩZ5�7Xۆ���[8����i����?�:N'i���9�d�nV!YҗJ6#TS�ڌ��.j��)~�\t@�?Y(P������Sg��='��#`+��5Eh�aV����$�7aA����*?A��uI(PP��ߊ���:��%�]Mϯzd�節7�����zz�v*����X�3�|�mMTe��gu�%Cb�ն��*N]�Kc�ca .�����^h
cJ�Qdqը��9�	�L��*!�wvl��@\6�7��u�D�bYciF�������>�m��g~�5`c�P�V��k�h�Ʈ����e���G'c�	�M�p]ʝ�~Ϫ �\���4��orW�gqѶ�~�7�<|�P �j(�����\�+�i���T$�ݒ�-����A�H<�q	��Wn\|yy�F�xf�����^�L�2��jAɶ��X�0�d��0좿��8'd��䑂%5.(����|�:���f����9"kxre�����2�̷���㷔+��%�^�f��aP^�i����e��O�i��#�s��^O�!��p쒜������u�4�7oA�4��f3��dM9J
#���Q�CH�O�!	��H���-��Z��e��	>f�}x��Ջ� ����L���.ؑB��
���0�>Y��x#"mb"��ZV��7�T�S�M%R0��i�M㲴n��}G�j�8B��գ��/jA)���SR�?+�@:�d��&abl)�N����Մ�SX:ڋ7�Z��
5/���-1�q�,=��}�8� Ϝ�ѧ���r����UF8E���n��4�k����̠��v޻���	���t�6�>ȑ�ݞp��N�iW/���ֹ��oa4�x>)�X���ɉ����&m7_�o�J��`�=�'�?Pel�}w��Ȅ �W�Q��w\���EK1�s'�"+]�Ͽ�k&6�;�Mɀ!."�O�Kؤ2
�qZ�p����ؙK[a�-h&��P� �pХ#=��er|�n�-r���b'56e��r�'�����ru���,�t��?�Ϩz�c�C?��m����J���Z#�&�����bo��/_����[�(�����&�ɂ6���n��I]!�{\K�se���E�[q�?��"�V��:[�f?�N�r\�z�03}��G�DF�\��D�{%��
Cou��x� �zw�@�dcgo\��̹wA�e��D7�Z�t��I7��y���
}�|jE9[�/�z�p���ϴqUc������+ދ�=w�L�k�4tC��Mkwl+������o~-�.�8�b5����e���Ȣ�]��M�y?h���4;S���2:�Ѱ�� �̥3�Ēt��f����F�7�}b�<c�Q���Q`:�JESuΙH�jڃ���G@��TE"%�>�8G4��J��P#��fq��ׯ�e��FD�>Y?��p�[Y�NU�����Dj��B�B?١$���������Ň���J���~f\�~[�������4�a����[�r��6�3p`l���ǒ�NƢfo!҉��L'l�b;��G|N#�m�ݒZ7Z�-�v���ה�Q[�QA��(� � �����憩�
Ox�:�ذc+���e���=�+�"�E�v�0�i^ZuVhw���a�����6D��Q:�f���{l�l�bo�>"M�i����흝&gW�L�������\��#r}�>y�D8���G�S������_~;V�bu/�d<�@T3�2���W+�&<��9H̥n*T,��vr���"�J�
�0�:X3��ǜ��QGGG������
ʹ|��K���2\�I��Ss��l�漩�M����\��Y֗��J����nJ}�tT�rpK�����M;9h�����g�r�/#l�-����T374;;[&��������,F�(4� �� \yc#���=�W�V����U�b{�KN��[4�T:L�+� +Z�����͛�2�c#�	Y.��'�����G�@j�f���BD��?��<�!:�pk��ݖ�NV%�
����HW�JU{�����-s�)������W2�gfV�w����Ag~S�g���!S��X`h%���w�v�^Pj�#Zdk~�,_���v����2����{����|���PF!?�?5uI ��}�E?Ϻ�1 �K?/(Th�*�gb�����]�0c�D���ؕ
s�7�[��M�(Mh�(x�"$�Ĥ2�/�/���(��`:H�o[fk�{VU �0���W�=��)z��h��sk���NmH�)�t���M�f����E��N`����Zg�pL�c%��W��4�9�b�����4��Y^��џ� YJHmDC0e��x�[*K�d�υ�X��7�yU s'�DN�%�?�(E����3�
��h��*4��b��b�B��4���'�F,.S�����"w=_A�n�ᙙ'f��@�����v�_I����ş!a�rI��B�.s��$��eh����}�#���h��6�|����5+��n�b$L�	#��C篽�z���|�9��9g�g�g���>1�ε��"n~3�Y�>��Y�y�"'f��#�hi��L9�.�P�S<P\r��3�aQjS|b.�t]bt�0���/�������q��s���@�|��sctc���ޯ������u�����	e��Sw�j{#{��׷ǀw;�|��L8���g���@�p��KVi�v�ijh'�M)ֶ�zS1zŁi*��N.H��LG,�X�R3#���+��>CJiz�oXD\*��mG�������V�N�5�`�'��%�?0{��
Pm�ߏ�[�q���9Cz^1�27dX*z�T�+�r�s�:��i��>�
������e0��V��h�s�N�M�����#f��0����`�*�B�]eC���_��%��B�-�Pu�4�~�$E��&1�4N�ed����Cޗ���Ca�<�P��s�l�N��=�W~[d[4Y�쾱�瑍�&��H̡\�?��?n� �/�b��=/��RLw�^���8>�e^o��n9h�(Mk����eMk�;Y��)�'A!���+gX=:omM�ʽS^�m[bS���u�WK�0���u�hC�E���]�8�����vH���Ɯ "��������]u�GF&	A��mXC�f��2E?*m�;c+�{{�q&q`��&�#��-���?q��F(U\ߙ$Ɓ	M���ny�ū��'*�5*_�xP�SYRY-E�?��)����0�l ���U�RP�����V�p[{���������]��(oi�^�l,���W�Vw4?��1J�Œ�0:>�|��˧��b����xuuu����;�������^�(͜}�b��tZ+��N�m;Wa�W
Kʌ�*"������a�ܫZ����
��Is���Q������2�g?�^1��h��z-��~Xi�������Cǔ:0��WK�����^x�^�ڢz1OFFn�X�#��5/ݦk#⎴�jO �v���S�	QvA�1-2NP�e��8���Է:��c�A$!,��}��^ay�MK|ն/w�rn���4����������!~�V��n��jՙ鷺6l���Pú�hW���;n:^tU�ljWH��?�AF�	kn�i����k	�:�����_v�/ˎ�,G�'�ˉ���Bk�w�WLD�d -?Lvz�Ҫ��<m�(ap��n�߿*�Γ�U���y�";υLy� �_��D0�.\���*��������}42�ԏuEut�-Wc��Xب�2� Y�"�s�V�R緭�_��;��KtQ����!�;Q��̰A��*�i����aXҝ��n��]�h=}��G�V�mz�׊?f��~���edK�ՂS�FMπ)<��w�3�!��Y@z5��Ħ��M)�2gd|��3����Zל�" �R���DEE��c�Bσ��m2�=�r{���V�7S"���n�=�H�2ʩd�����g,sw9�,��}���v���m^
�gΪK����ܵ�6�u��)ӓF���V�t����p82K)&|�W'����{w}C�R����G�� �$�x����]qV�����̒2m����T�ԤW>�>�B�T�mK>�%yL!D`�ć���cp�[H�8CO�Ͻ�@]�ɹ��HNBs�U�(��nXQ�^��:UbS�i�6"���S(k?q�����B"�4uuu�<(>�K� 6zfN��1xi񿑑���{�KA���Ox<���~��~��̭�gI�tmr	�K��^����D6;w,��Z��(��R%��(3Z�ܶS��/"Kd�#s�{:!C�~�Y�*�t�4�f�(k?��ÌR4���3_��w��K�8I�v�E��۽6���[��R��xHV�q�>|����F�{�<9eB��v��L���M�J�+�G��+�$������n+�&�e ���^ �e)���|K������F��B���j�y{&���;��b�
jP4����3U+Kߚ�+�ac�G�N��Ϳf(¿BVk{�}'��u'��D��Mc�2<�S�cg%@��{~�I$�)0�T�]����	D��O��)�Y��@�r�"��P����3��.�����Ş������r�:�%0���Ҫ�_ih6�ǝz�iL,����,��rs��d��X����;��oy�:�L4 �Y���9CcGJ�DoK2�&�`2Oco�+�-����Hw��%,Z��D�!��K��q�~aʗ(z�^F�W~@��KSc����{�C܂����4Xο�Uqፋ��Ec�<��������^����,9e�G\���k׳�ȩ]kl*e�˧
Y>���D>�ql��cO�hmi��)z[�� ˎ5ʣ�hk'�~��,�W��~�����m2�]{2z�(ьy����膄�P�I	ϜL"q�Lƪ�,�<z����'{��1�^<G��Mi�c��
B���y���	�{�Vfn�<r��>�㯱�L�ԑ�}��s%�ȶ�Y�|�y���n �:ַ���'�I����!����/��ؒ����o�_����4z7��}�*�d��÷5&(���k<%���{4M|ѵ��� ���K�`�B��,����ˋp����k��=����QL�4�d�a�����Ewf�L@���T��ؓk[�+��[ʽ��'�J�h���4V{{{V��ܫ\y*�'�b�"����2��sb�AwG���Y�CJ瞤���R0c_�קKt�x}�<�yX!^Y<�9e�n���4-$���充��}	F�%��������J�ˍ�KcA��߁��9}؈�s%�=1�|�/�=�J5��T#2�}:��Bsణ4'.��Z����?\��~�ChxLJ״�56�%u��4�����/u?�?7f�Qv�x*�dSFy�����^P�����L�����\���χ���%���#@�pr`ڙ*���a��~	,ű�nW1��\c�1~�����}Iw17F�'a:�+��2�ZߵN4Ba?�;�&���E޽�|���QE�����vkN�|��qM�x@����e�U�dT"e�hf�K��~��0��kK�GK����<<	�"q������5��c�΁bƙ�wE>��Q����:@�+0�dvψ7VWGB��\ϻ��li~Y��v=�r���$m����Y#nz&u),��#��Tg�T��j�dv(�ڴq��cǾ8���1�*/l���R�����!��A� ��EK��. �P�h�jj�2��7d���zΎxIlಙ������K�>����|�������ݳv*��(< �ܩnͩ���^�.�yt�<(�f�������x�3�75wۙ��b�,4�������}����Ty�B��:����=�2�z/����I8��kh�DWť��#�߱�@���Y�]rp�/">��i�YA�ݱp"0_����/��!�<��+�<����6[��Ɛp�3 �6���Yb��G|�1����i�M�f*�ǻݛWxKx������b�646��
ۓ��a�C`=�XD�=�����.�1�S�՚���r�7�㻾X�@�Y}X�>�D�u#��,	�ݷ"~jQ�����Ȇ^F��.��1B�I︒��f%�Ib�e3��Q���/C�o(�����n8��l�j6�lGwS�9D]������KE�i�ˤ���j�a���Ws��9Dd��44h� M�x��d�Ω��4�y&p���=)�׫ ����^����������ͯuM~_������E[�ު1�K����39hpm+���r�6����hl��Ş��@p���R�'�A��>b"����dɚ��0�-�5N&��N����ȥ�u�˷UL ̞U��l������E�:0����Ϲ ;���d^�٠�3ݙ@:���a��#5֏���¨kפ��g������)�;q8�+0�7aIOߟ}G�6` �$�������z^"���j+��XӎCp"T 2��WC�s��/���E>�	Ѡv}��H$�*]#^��$4m(��Q௏Q�����yW�'�!Zy$_ tDҪrx�)�c�Db�� k_!�/� �HK��1记ng>Gի ����0r��?PK   �yDY���  �  /   images/5d57974f-fced-4f10-a93b-7d150e366d9f.png��ePN��)�
�J!��"-<�;��
���-����P
�)�ZH���^�yy�y?<����ٛ�ٽ�۽�E����```+�Kk<i�')�>�~$�:O
�I^�����+Ϻ��4���dt�4-�<�]�1<==�Y;غ�;��st��9��``І(HKhy��y'�n������z5@���I*��},4"H��=[�俜��dVM��������z,�����L�	����S����q[pp�_Et�fe���9���y�я--�V�X.V.�]�����Oq �AA����;���%f0w���j����GǇ��E��0�?���RY�u8� ׫1�MMi����������X���M"���
8��:�����w(OQQ^Nz���V��N�A}}}�y��A_!m0����E� �����%e���#��CB{4R��/��}F�
�f}� ��%5EE�����=q�P�E��W">�ĵs�D���iuuu�����OGk�
��D�����Y���&lW���s��>ͬYŁ0V�/��"��I��	{�'�
���H(���o*�^�I�q�QQQ�s\U�I<����
S#�5c�7A�����ϯ$'���;�B��>��5�ׇRA����&�~@����2c���R��6=Z$�"�y��A�r�����^�߉��IJ	*�0	ua��JХt ��/ő8�1�4B�M����l30l&�^�w�ϝ��19�٫��!!!��c(&fg��2\��f`
�llE%%�Ǔ�Xw��1�������?jyB��Ow??1=������I8\���+ɸ6�_����9b��)�:	i�
�\F�c��e55�[�$�� ��O���Դ�����MM����q%E�B���!�Q&���<|��ں��(��輄.��ʪ��e�[~Қ����Q�;��*���B�Fe�����ܓ��[.?2��i�ج��3㹵��Ժ����%���ե��xbA�ֆ�)�js4�������D3�&S�p82R�;���w����6��C{`ek;6)P�![�%�а�i�������9����_�5A�DIu-����wpI�@��2+a�����h�l���a�%�\� �G俵^%ooo�R��Ut�%����)1L�Ǡ����� �=z��G+�Y%��t����T�hSJj`�����}�v���&�o������b��y1�r)p�/�T"�l�7]�B�������(Tl���E����!50��H���|R�-�8�����`9%e'�l��s�����C���� ���=��Do��K��M��+���J����`C9W`��כ9���7�{�K����t^���3=[QV������rۜ��%	~��}�q�b�SJg�]p x��L���l�BTש�I�'z�>����Ӓ0�]��'��A��z}R.vG��Y��<56�6�������Q�R��*+��#sgý���?�D��J�����v����2�~8�fȟ��J�^�Oє�~a�Iǰ�s�^[��kfs�<y�T�C5!K�'˽�Mv���%ǷH���q#�pۭ愅�#ua��O�n� �ډ�����N H�����i�QD����6���h]�<����¤��w�zv�"�n�}��X��o$�DI1�muZ	�#��b����sC��*�gcs�a>	c �a�ɤU��YH���[u�p#yP��q�sr����*��w��k���24�@^
%?̕�dX�����!E���8z���:�d.�TS��%�M29U��֐�AM(���(3E%p�W�2��V&v�[0X� ��m���[� Oێ� �����������!���X+^?~�BI��01Sxt��s����G�:�;/̉K�p����f�_��	����>���:Щ�+1�-+�2	Lq��@�aD8� ���P[B��l���h��R�)|c���<�����B�l�bˊ���(���_�e=��bE>�L��B�%e�`���
y}�Mb>�+H6̠J�u��ZE����/c�+f�l�a�#��g�~d2��
�hl¢����ɐP[��43�K����A�~��)�^$�~0���oss߈AҐ�k0+����j��S��W|�V����Y�$�/�g�!���E��0&2�������+�"k�6yZ	��ѫ������_?��'K��:^��~C��;e��J�D��|��Z&�]���(l�@;��Ӧ����t���/�.�\·p�@VϫD-��?���n���vHb`v��X��'�,[���|�U|�Ö-;~&���N���p�g?q(?��=H�YP��f���Eka������yF�.�_.��N�E�o��:�`�T";Ló�w	�}�5��k��F��x��hz�ߝY�7D_��{u`4EMJ%d���eXEepbz��Ds\����
�oJ�=BG�~�AA���=���l�ծ��?J� �;���B�T���<���G���8����ma�R��B my�-�J������U�Z��[\�f���Y|e?��_�F�U�H�o���oz�+j�����WX9���%�:	��$#�A��))~��dϢp�����5��/d�C��P*�:�}��oV���sL�Nc�VWèf�%Dom��7�E��E�˾�9ZG�Ӹ[�_;KQB���$�O:�9Y�<�W���S�o�3�P�<��iSuG�O\�(o/�c����-�;T%W md1MU�⾚L��%p��g:h΢uXcI��o&���O$�.D��t�2*�:��/P��x �CJV�N#���F���y�mb�r�x����3v����W}W0~�#��<�Wi4��P��ǳ2$�"ĝ"4�������\(�������ҝ���A ���ښ��%+�3!4��Q:�ۉ�-`�S���G�k���A �^����n�R�����ܘl�װ����S��2�W�\�+g�\��ɾ�I�� .���l:^����C�f�EE�|=�ϫP��.ϴ����bɝ�:} ������{ggK&�&�h��n������4�(	N����+%���%���i��7ۙ�RL��	�1�w����-����Kf#ǟ�'�i��J����K�iǓ��\� ��ծ���l({_�1ss}����!:>�9.ڕ�A��~�����\4xd]�DIS��ڙm���'P�\�T[��6�z��o{�J���u���P{���Mv;ԫ�F9N�6�$�#���J�DI�������y!!K?��/e�픥��°P�5�t:�P9Om{���@,��������)�D��·�oiچ�-B�Hk�g�{QPHTfn���4\6N�;"�����ʚ��cTy�Em�t�q{h,��f ���lllB�q���C�PV�Y��X䃄��3P���׉LbiŠ�C�߈]u$��CE���K��S<�ZҨ���X9��q��Դ*��>�
ƜK�ΡU����4�Cv*���U����M +��BQ(�y�&a�t�UC���#���P#3�$�D��)q�H��$"����<��
D;6;�A��af�Uм��ikC�b"@��5�Z�g�	���)�Ǔ%۞Ue��@��e~p��K~�ߛ��L�-�s�x�d4Bű�K�_?�F.=kwK�2��Hn_�*q���O��K�o�������I�ef�|�&���|���x6�U���n�Y��A��xK��g᪩Y�%�TՒ��qi5R�^����aMYރR.#���v�~}�?~�����Z���)Zp�BQ�,�~qY�#�W���^;^���t�L��0�Ȋ��ddVQSYv��<�xN�*o�y"�)���`�;3'��g����2�*vJȨ�^`��O<��p���f<��05� �d���=m��3�a�Q?=�̈́7G�&�J 7hv(�@V������Щ|ѦYQ�[�d�.��X.ޣ4ە��$#������I�d��!0���kqQ��C��M����#gzb9R^:�R�f\���u_@;/�MNKdlz����F?}���pe���<�D�t���O^��g���&AAYAu"{�9Ec��iRϲ�d/{�}ׄ
Ҹ�;���~�(%iC��:x�<Q��㿽�ɀ��i��>}��W$tB�W=��c�3i��f�n��>..nx _�5�/M�b�3�3�ua3Sg~z�z����]A�~g@�W��.O�QBHHV��w�4/x�R�;Ҽ���G�x}33��X��Z�89��Z���͝oy,�x}FٟH��A�?к6�:܈�3�P�r��O-@��ݞ�F~*��8�*��#$<VXcQjٰ��L�Rz��Z>�����d�W0{�|V�uw}�x���:�M�A��A�O�s��P�U���p��S�a9j;��w����O����<�B i����\�ʥ����ˊ���v�q���Ӊ�!L���M��R��A��Pz$.�D���������Kψ�߀yO_Q����K��M%���z�+���<L�^�]�����<Ԗ�Xo�����ǩ�C!$D��Th1�Zڅ�@������2���qc�Õv�tܒC�Q	�[�g�q���Ka������7S�r�h��vm�#b�7ם�q��ؤ�O9�Z���P+����>�/v���.Q�!��9
�<��FM�0�l�Q��LҀ�h��˝��D�)�fw����DQR7+On�ri%)�3�a�Œ�<���̮ʏo~�R�1�6}5FBdI@�(ݛ1��L�G�q����N�A}]H��Z!R2'�o�1�v.���.zw�͢BP�9
�|��"F��o>�W';K��1֎_��9 �32�,r�i$�W��1�_I�9���>z.�NZ��ml\�۞C�ט[�{^�5g���ʙ����WNm3爛�����'����A�c�2&�q�������KM���f,K{b��u5f�f;(v�C��1~9L��\�-ӟ@��`��%�,Rx�u�l�#1.^Y�"^�?E��v��m�����������)�F�NS�����E�A�0�8r
?|yn%m u���W���t<���>����)���ݴN1GQd(�{������@`V�e��� ���EhXx���pR%�`3p��R4���u�M�ƌ���f1N�_���n9T�����"ǡ�|�~m���w�Y����.hvzA�MhL�[�W+:�~�^���ť��K�`6�sLL�ū=�z~<!a!{�sL����+%���Z��F�mYU�{�jC��l=����<�gbP1�E�GI[�o�ER�ߒ,���*�e_L2�bi�t�I$��b��]olƼ�ju��T�t�L�~UGo\}Y�oъ�6_����gU����=��A��}H�־���F�&���i�ݯ�&��(tiH�d�X�U�!H�ТR4t��mi���ܠ� 9�u~;���\���n��t�{���	Ҫ�k����R�#�
��y�q�b-�3��e"��o�:��es�_�� ݍ�:&�Y�>�a��wB�ls�����
V��?�e n��L�L˛2o1}�F��J_��[�''<���pYOffЛ�j�G�u,�� .�����NnYV�5�w��	�'FV�d�$X޲�nV֔���`jֲW��\J��X��tE��hh�3P�m�N
�A-?X���nܳ�R��?U^�WU�m2.���S
&���"����{>j���;QP�|��F�����2>�E���M��v��
�ohؽ�99\ S0��q�1�*�m䕞��}�?*/��.�]=6����#A��%�V���v��ư�J၃��>tJ��9[S��=���)S"���a	J�o��!�)�If�Z��9z��@Sg7���Dfڀ����������ť�=�"KX]-�ȑ<��Z�N�p>��7�y�l)��/��|����?�}a��Ŵ����[ ���"��E)hOVm�`z#�RVq9wpaط�+�Y��*}��� �=���&)�i�J�P�����+��~]�eܤQ��t�wxx8� ��-�L�[Y7W�<�q���G��kN�QR��cc�Z�Ϯ�}�Ĵ�f]؂֡��7�FP��9�GyW�ŬmYa�V���Accrw���~�S����c�[��PX�����Zg=$�\�ʦ��^�h�w�t5��hS}�T�1H�@ ��4v�RQQ�p-�<�D�_�1&�C^Tf��{���jX�x*sߺF-����n��9e��i��/s���
p1���c
E�>���5G۰��R��,��w������8���������!R��P��R��N���W�T&�j lx���&�* 3��B%�&r�����7+�Q���xev�;��+��w���k��c��G�u|�\�2�6��á�c�Z�QKCS�s�ݴ��;7�#�"7��1����v���.À���Z��y4<�/��>��l=!�n-E�ǒs�
��Ε�INN��*�[����v}��kuu�t�zO�,	������𜆻�0�8KJ�����1�g�w�;/���~�s�\L`��
rx�U�7�Z'�'_1����B��ll��nF�g�'Q�`)�4'E�5*r	�Ͻ�m�倵�*���~E�	{v��F��:�W��!����^�V�۝����KD�\ӽ�C�������;	b�;�e��"����L�C\z�c*Zhä����y�zm-�u�]�<�	�[�H��5��_�D״,��	�w����kˡԡ�]���ᇼ�_2ٯt�5�E@�0c~���_1�%��,l�̮�'�����h�)E�i������뚺�]^K�)��zHG�>'�7o(+m��R� �8hI��Oz!�0�������,��b�7��&�Ҋ�,�އ�<[��+rj�%o��<V��q`�g`_tT�׃z��U��wU�{2i�����啷� ������C�I������C�Lg�Q������S���S9�_'�Q��*W-�����|�\��`�A _���� �*]-i� PK   �x�X��/F��  ��  /   images/8278d802-2c3e-4ab9-9a04-8028f624633c.png ;@Ŀ�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi� @�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:��� @俉��N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0���7/�Щf�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK   �x�X�ة� � /   images/8d398a91-1a51-4737-8347-b2d4588b3940.png4Zct]]�Mnl'76۶��F�ƶm�qc�qc�N�_�o���>?�^{,̵�<gG*+J!������!�H��~�a``���_OF �̯�EUJ�f���LF\D����/�������zje ��} �,"
^K�v6:
6�q3:* �6�@|P��FED8a�K�AM鵷y
6�9�k�q˓��s4.�����{b�7�sR�������r�xm����	5���x=�$	VI��\Ҳ��L��6E����ZܘTIy�c��4n����bO�������'z�<�Q�w�ڹ�[�@��p���UܧJd��ʑ�T&���Ϝ�F�\�|��Q�Ώ�o��������M���NIg~�5-K�??�-����;��C�Y ʥ�W�8����xڋ��G�K)��Sq�U:	RBt�O���eP.��rΧ��3��nN�~�]�%���L����9g9~�@�a��z�Z,�'���[��"@�aW(5!��X���d����z�-3�c6�,��T������P+�);�0Bg��|a1�_`�@~���b����'�D<M��V 9����-��\��:�	Јh
Y�P�}��d��ƭ�;n�+[�Y�{��9�y8���Z�������^��lG�k�I���o�]W[N!p�]/�Ur>���I���,	� ��9v��/�^;)F� 1���u3�UT�_���#����������ڟ\��ܫ�8����͑�v�����{Mw�	�ם�㳹�qu�c�)`e��/6:Q���/zɮ���� L�p�<���,ב��v���G���ڹ!��G�'q����Z%Y��1�]��ޕ�r?�)��t-&��]�5���� r@��h�y)v�;�?r`�D46��U?�F��?"��hʧɲ�gl����bŲ������O� _� �ƣ�n�1�5��T�<���u����d�Bm��JGq5tj��Xl>�}3s ���ےB��<5O�e���HS�y?�>�-nw�n�2�S��~R�q���k��k�$	UT���n|�{;��5;�y��Ñg�
����,r�vc�ߠ�Cvχ��1�����ٸ=@Iĝ��Pb�.&a	ݫ�&���|��|�����6���P ��i����u04R��pM;��.*d"�T���b[�4Be�\`�G>���z��̓�����y~�:�h�Ϋ̅*�-��􄒈�S�u�Ɛ Ih[T�U%�w�+�'{~5p�?|��wv��Y��*�y�8���5�p�j�k��&x�i1�I'!"�C#��Q+M}�/�
Լ��js����a#3�]�+*i�4c%���
dLɱ�ط���[��Ϲ�QQ�z	��+w?�w�xyt-�if��ǆ�	�&CM2�Y�D�Z@�:�k+Z�F`�=�Y��Ώ��]�,�ޘj:,T.DVy���7���!AE=��u�D�&;���A������c����H�6L�T����f������}&�5:|��5��FF.����7z"c#�Q�vvfQ�}����W�g�"��q+�ϲ���[c������$.#��x��ސ���S6�jA�Qx	�@�rG"��R��{���S�U���x`���x���[�R��N�Qw�\�5Z�L�h>4
���/�%�x�7V�u� �,˝SFe���Å��� ���v���!|�-.�oE���?9]Պse� �\��찾�db�`̢|�M�A$�s�?O�	�gw���%�y��u�ʵ�s�ړ�1G/�f��?�q߮�#�OР����2�حg3V�!��`ȳ����tr*I+Hǰ��s�M��̮K�;8;f��:��u?��j^�q�F���'N-".���Z�o�`]|���s�Ƀ�F҄a�I�67��6d*�0
���r���5zT1�c&��~�B!O����L�`9h�SV�9'�T�<~��R��TEEERο)%ï�,
�������j�����j6���z�-lgK"�ڢ�"��n0��MV*�e�~/��yX\&����[���f��fQLLLL�Mr� mM� M��U�|����#O��8���~�E���{,ZbF�v���J�a��h9��6� )���v�X�b��w�!L�u?���Jn>]"��;���2���b�N�"����\#��w�:�M��?S��?�ɿl5��|�����.����cL��?b���D�E������E<�:��r{���,��H���50��^�XMC�����d�	�_#�����A���6a8r�Q��o�;ڒ�������l�ۆZ֖:p5^ȯ�\����Q8�az�0�+�c{m4��[æg�|W��JYx�M_�.�j����s .�h5XK{��&��!�A��l�{P�Q�'@D���ڟ�y��ّ��|������q��n�d���c���#����i��0�9ԅM��n�-NI:�d$I���ta��̽���$6�<F����@Ny&�=�D���f�������z\��'@�&�Bl�c�RC)�h�����;t4T��]�1 ��6�4 
���P%&5:�L�%x�٩}�UUltD�+]�&�9�7��	I��e���*g��kb�4�'�=N-_1�/�Iqt���)��B�7/[�T�/���N�����ҭ����or�u;�Hs��p1	���&��t[k���F���G?�K���Mi;u(2[<�zg�T+c���*�4�z���J���*TԶ_��Y���^��=��D��1@����NMK
V���]S���,u&��qÅ�^�4��m?M�5�չ����&�|��O�>@�r�����72��]k��y�#�����+�W���&.�O�����,C�8o�D��Y*A�ê>t�Y8G��^�B���N�Iؿ+pq*���Dw���2��aH�hhp��9�ξQE�����>�|B��>����>���[�ya�����;84�lM����$����J%}��$-
+Ga!_��@wI^��IVlF�$"W8�Q$�I�}��pJw�M!��?�YU]a�/������W_8��苙���ҰP�N�6/z�he�������(�*�%�"Nv��R�����@�&��݄��Q�Y}��.ܗIʌ0��}�����W�x����#o���X0-�>����F�~��;�8"P<KV�)�"I4E7	�
��+4�r �M���TBr5�g͎���U����Q�Y&�g�-�:�3�9���K�^�4,p"��*6�J2[�0��e""-�!&^�\��6�� �eb��r�Y@�\��l��C���}a5"�Z�ʎaE@�KL��M �������F�t2�:�pA{����pRI0�$�h$�Y �Kd�K쥮�������DI��AQN�T�v���ɜ�R��׀H�M��/�PW�זv��D�]�Ѱ��,�+���I��T��u�):��de=�h�H��}�(���qK�h�!���w)��Io�C����s#���q+l���$	�~@�0�r�nt��{O��6�S�L�^���"��<�Vj�����F���<|�^ry��p����|��P�0;�1��*6�]��Nl`���Ѐ2ҝ���L��'.��B���oo0�dk��l���+p��m��d|	�ߢ���n��-/����=����?���W�����O���!cn��1��~�nڰ[M�@ 6�<\l��U�~�ol�D-��cZ-?e(ANaŒ8G���w^nmK,?֨����z^/��V����.`���VZmǦ�Ă�k-�d��g"�uڄ�������jLH���� �<�|^W�~R���V|�H��+��)�8,L߫v����t�*�o90h���M�G�/nޣX�7�;'��n�{D�n���F����9�A���ōy�n剌������o��]���3�O]+S׺�U5����}��G���2·�n�н6�`F�o��4m6K�l�
U��	��!~����%C��L�@I0��ﴸ@�-4���l�WO�b�����>#�p1	l�7�T�aH߆Au��}0�	W�-���N��%SB]l��6].g�}o��j�+���5-�s���^,��,�"K��{ c,�Nb��[�y���+4��~���h��Ԋv���#[��D����21$�n����8c�5�Q�ѥ������Ui�U��]�����g��3�` ��bEt�u��I����鶱����j��r�뽲��l�]|ɸ�8��4&]�s��:����_���/�yT�;��x9��!�0ZK��b���/�'�pEma�܁�E���y��Q���4)�����'��`�S<!_K�r�iz��G#��d�j[�������XG�p��l��e��|-�.�a�>��4�Ð�vޝ��_�o�������f�z۲�	��@���J��Zˏ�ƛ-�S}����\O�)�^��ndM�&��&믺��� ���.`�nz2t=�+�E��e��n��[{=.���5�wd�3�K�������»�4H�ۮ�X���1�:5t. �Ǡ�ş�m5Lgԟ1��`Iк�����p>���x� ����G�����^���d3��zI� �)���x��*g(Ģ�� ��"��&k������􆾶2u;et_r���8�D{7Ϸtl|(6���0CU��$�X��qfj��B,Ds���{<�I|a���\(&���4�=�j&�֗^6b����v3��u=�o���#���]d�1�������e8�Fa _���/I�wO��8�S�ߺ��?�_�Ϫ�l��Y�à@�_�m�K?�y8��yd�}��`ID���*�ϗg����n���B�jΙ�bD�����Z��R���)�k�*4 ʹ�>Ë� �$�S�4���tCL�5���y�S���ƺʌ/ �db���j��u[:�#��{���������s�q�[��b����R�3���܍����" �	��{)8�bp����
nr���������l*�*�h��`�;~�nX��o�f*�����AI��Q����.�i9?���oK��7�O
�Lh$���/;��q������:���>����zpF8��=�xC��{���uu0p6�|JIIa]�S��9S��X����r����,�H�Eҭ��0���Y�=� ���`���B��82�����7��	�|n���{kT<�N��3��l�PŻc��'��p�Dd�7%P�,G��~o�/����7�t��C$��:i�K�;<��
s����cw��26�h�ӵ�ï^e�l�Q��)����xG%����^
׫+9��A����8X>РA��7��R��8�������1��䴖���B�7k�]�Ͷ�-Xc��V�`W����/\r���z.{�_jGC|1^0��y�����9�eD��${!�Kat?���׹PB��0Vz�����t3���LB�s6R����;���o�?$��[��T�h�������E�ea���L�����p�\*.ǉ#�a��VM*�34@d���
GE3�H�&�mk�G�sL1�M}���8��"��G@0������C�Rʋ�n�_轤���~x�s�a1^gꭾ�^9���f�U̅���K���D�L�ewI9�k�;�e.�~���9^��#t�]��0ŷ^�
��������K�/L�455m��K���2��ٽ�����>�"i�<��nd�A�r�p���YXƕ��z�N���:���TR������V�o�H��|����D!<��Т �p�}�	����M�4�^����V�>�ߟnl�����w���+��5	�FD<֫���ȗZ�˵2�/������7�,ty����������� �ǐ4�d������Xu��ٖcBFΦ4�p��W�d=�+��={�����R_a���[g,���L��Mжo��(�6&�#JƼ]����i���b���_��-������@a�"��r$՛�Q}Ѱ������V��/>"dڶ6V����f��d��`csZY�ŶrA��5����yt����&�!��c�N|*�)#E�~6Q-�2DI���ݛ��j5b܂��H�.��q�1gLR���0�;/���ɀL���"�?,c�W�|� j��b�%o���W<��?�:.q��=n�~�� c*�r�D�q,�_�u�V8UֿX!*�؄;�7������U!��l:r[`�V�C�l�o�)\�K)��0�v�wi�y��	�Yv�]�}y���i@��d*:�ʐI͕.sb�#�h���%X�B՘�O�Ӝ��:�����G�)�|1,'�U�8�����N��:Z�$�����*N�A�i�C���*�gZb���C���@4���

�}f"��<��]��{���ֵF_AC=�H��ߚ�*z��(���[m�m�C���������9��d|��}��v��`bη]�L8j�s?��uy������ר��Ld�3�X���|N}���ÝLw�������p��siA@4��{�g�H��M׵�,l.�N��Ơ��[�7]��=)Sʯ��D�]�J5z=#E���b9��r����<%fZ)dF`��d�Z�C{��{�m/�p7�H)y��N �uW:��1֞@)�٥��z�"�����7��\�_�3l��w��"t��dG��ZK|(R�N��%%!9r%PA����-��������6�к��h���E����]UV�o>2Af,��p���."#`h����l���"�y��@S��*j��<��e�)�8��&Ȕ/R�{���jCmOG����?
�II{_ܜk&(�k*������`jh�iXG���l,��M�w�$�O���o��ttx��u>'8�M�����~�/��[y�6��v�E���&��t�f�����9F/����Z��{kD�~�f�JJ%��!��f	��=U���q����Xr@=���+�9��\�U�Lq�٨/h�+�G�~S��%��$�����.~U���X��,�)Q��$��UV��5��[f���쮐�-Z)�d�I���P��M���r;s���lv:��F��9,V�j�ֻ��]�������{Nl�D7e��{=_�F�y�3Z��޺�2Ԯ��X�9%�xT�մ9��tj��vE�$��~�wBq�\,6�5x�a8+bw��y�*�_��<M�� �X,'s$���;N=$�A`�W!鯁md� W}k!�g���ʑ�U�
�eC5+.R�8����T�'��ð��5��}h~V[x&`�:�i��>��e	x?���~챹��3r�O�"i2���`d'ʈ�^^��������a�1���f�[������n�OV�lۇ�0$|�p���T��/<'͑�2�w���Onfi���[w�سJZcG^
�#��>^B��z��'^K5����לG�RB���;#��21���/I���j��F
�y��|_�������s'�k�{�6 �Q��Y(�H(`����,LZ��4��J�1��?����s�^Y�+=��G���D��m�у�Q�Z`N:�R�5[��	zaT��+T�2G�S�� X�E�#�8���Y*�J�ac�
����8���G�a|����y~��K���T%h�#Ho{�ER�|�w��bL/��������9��h�(f��%� ��	��9Ŗ?�������6�?��-s�L2�E��f�	>�r��1�p��A�� ���	�j��ʼ�Ȼd��p�>��\��ǈ^�\}e�A���g/��/��~~���f���]a�=�-���	�1�87�x��p�a�E��~F4q� ����+C��_���#/�3qD�ԁH^��L�C��s��>���.{O�}�[9mJ�/��f�z'��떬�.aR�eh�AOD��by��αyp��(��
�S���u����_���'�2]\����l�*�>o���{�B&�z�b�ΜeBn�{�l�o����+���#~N�р�9�7�Oq��#�cLK��`Ez�U
H���'�"y�JcddtT��{�4t����0���Ip�"��O�_�'S)Z	�=uf1D��.�+���)�r����
	w�G*����*g�T�tw��x\T�rG	�Q(6�$�m�
�|zeT�����C!����`_�0��pN$��"�@>O�>��T��屼���T̘e�~���&����袂횰�Swn� �����K{y�n�%tlK�U��n8�����u�^�<>�-0{�!�!Nn��+�{m�g�S&U���k'|�����m�!��\1:g�LC�I�����5��
O�X�w4�F7�Z�]�C�|�[�� >jp	��,�Ң��Dh>ѿy|�@�k_:�F�Oy/�^?����8]��><C�oA=?nQ�����}	j"4������z��>7�
�ys�Q�+�I{w�������n~��z�3�}�L���M!t��h.1�?��������ƿ�n�������]�p��X���W�H=����u��2U��<��u�3L��ks4V0���+���Ԛ�'��f����۴T���h<��[e�}�������p����Ȥ��6>W��C^��ԑ�^�`�p�Ç��c�,"�U����ް�С}�XчըT��B�s�;`������=�c��ӧ��zi'�0"h9f�;��{�L�6]�U�����}Œ����?������F�<���Q(�F_ߎ �
�o(�<��-�>[aXV=�34�p���BFͣ!��Rs�\o����Z��z��zR�q3�}˿[;�[��)�����k0�M�l҇A�����{����t�o��g�jH�����N�m�[xN\��f�-�_�w�]��A�WN*u���L�e��Ó�r"O�9�[K��y?�k�FjK!�g�ѿ}��-5Ԧ�_�p@�����ݭ�t}���!3�ϼvk��B�8��F������Gb����U�a���w�����رR��},��'8�{��P5#�ft���5�:9¾��x� ��x��P�\q�����"Z6��F�;�R��n���{0�57�$�Ӟr�+��4Ň�y��`�d4��� �D�4�L"jz�H\dus�߼�P�<
�c����D�6�=����<t�D�a��L*���x�2W_����J}u�Ο	kab����4b�R�{�����z�!���`�}�K���ߜ+�3qR��UmE����H�EZ@OӞOe󀽚�R�e{�0"2�ze��*�K"4�j��x��|����,��5x�8C��"�����Qnu�]���h&6�U��m�
<^�vn�U��6�Q5��������	�f����	}al#��QM����f����M�)-�&j�B<�P�=�,���G;{#��:�HO�;��"ϯ�=���Ѡ:����Cϙ��ُFaI�)��t��Ym�qj~<���{�ӽ��y3���B�p�mk�G%z.5����!=$$,b�-d��e�����,�G�?=����I*�*`�*�*����J� mUs�.�@��x.���63;7$
z��*^�)��65��Nl:�j��a��m��rPJ;�svɆ@�9��U#�C��X���ڢ�m�������zG�+(���G� :4zM/Z�q[�i�W(ɡ"�ߙa�B����g6ח���C���H���b,��X���$�:��~�`���)[0���}�IA�H�{�d�27�VyybYp�°�_K#G��9	X�4�n�b��vgj=�EAMy#![�~�ZV��HJ%	H�"���.FMHv��;=e'Nő@o�x4�"JI��Y[E����Rp�z�E��(���J���]��H��T�l��NC�ҊZ�}��o�U��t�j`�k���s/��1Nd{O"��弧�J�y���޾�>*�W0�n��Y[re:8J�i���Kۻ1nI�׫�v�S]��uR��Іղ������[[/��OEU��ʰ[�FƧ"�D��P���*s�D[��B�l���}	g8��&E��� F߬�S���} �9�U¤F�����d��"D6:.���	0]�<|q�NZW�8�:���@�Ӑ �>kҶ�I�!s�o�8�^E�}��T��V��N>D����l��%�%��\�SP�(��y"P����u��d �g�+��o��(��|��A��WV�ڰ᷃�H�#1�q�$*/�"&��߾��d�>� ex�w�+jm�V������h�s���S��Cb��"��aA�v�,�ʒ�&�Q�f�K�Z���r���eW,{[,�&� �L��tkts���u2�H�l��'a^"���O�e$bh�y��z����#�r���%v�����J�sLFC� �+�|��98(?H���u�\B.�����N���+1I��_��&��A�6R�K�ʨ}`i����d���N�"D�uL�2��023�Z�a�h���=�B�iF��������� �fy����l>�ro7����h�:O��}{���>�q,v'��F�t��p�������,Y:�!c��Yga�tM�~6Y{ڌdF��j?�������z`֒�s�n`�5j.G�"�G���@>�Ó��KF:�J��u�f4���ϡ�F�>�]�v���Š�8�#� u���\��჉��q_r,bD&�v&7��.6�� B���.�e�N���g�'�<� �;O��%�qL��⟞t�-9��=�+X�n��pI�'��"1+�!��RS �oy�	�k�ޝ�ߝFs)�f
x;eo�QWw��Bq����C�!��^d|��b�*6�T���]◦T�KG�\`A�_�d[������,*�ތ)��-̒f��n�n��$�L#T�,�H{CK�O�- �P5�iE`�ᬾ
�TP��O�������n���G�(��
qIǱ��H�wC��_�;ϐE�4		�;[�9�˝'���+[��x����Xf�D���y�5�Tc�GrX��a�d�ϑ1>�z8����#�rH����М=|�̦ˇ_���� ��9Jħټ~?�Ġq��3D�-�өfbp�}�A���:P��i�=�v��\	~\�����p7���b$:��d�[箷 �%ʐ�ܮ��3]0�K����H�ĕ}{��Ps�P�Kn��2?df1�3����шT��
Z��w|3L!�X u�7���x��e�EN��T��9�Ŵ����AH:		�Ce�F{�������;�<�A��J�v�Y�\���n�|�+�׺�}	�.!�̇ëἳ��.E0��$A���'�_Pa�2ܭg��?>�
�й�i�ڻY�X�42��&}3�VDZ11�h

K,�8�CE������~5�`:n�o�$Cdj�-���3�	�!���Ա�/�C�z�z(`�d8��(Ig%���@jm�U�a<�;�0` 3�Ϡ5>QT˷n�a#h�S'� �Y�(�I���xKF�ЪX.u��*����̤@$��+(�K� ܵ�:��S�f0��!��t��p&�\���8���-��[hB�^�n���dC�(�\M3��l�FX�\3 ,5���*�2�;Nj,���p�ߑ���?��}�;�缀�f��,&�"��5 �M<l[�pΣ���Xب����E5����u��GΝ$YL��6��@���W�ʍ���s$5��NP�eޏ�ȅ��Q���Ytϟ �HN���o�>'��<�i:���d��?u4�`u���ko#) Ϝ��ʨw�n��´	��������#����CB�ӳ$BpH��uPW�0<h��t"��­�����,ǒ=��Q'�Ht��ۀ
J %,pY´t	����p�0#L��x��3�c��g\�|U�V�	lV��)�WD���L}<��0��#FƟj�R%�e&XmH%��U~�����s��kk�p7�ª�B���7䂄���A��T7;��HO �$K�<�*��d az�=d��چ;�E@�Re��܄�ǺbE�`%%�s�Cf�;�- d�
��a��<��G�3��;	B�4�-D���	��j�rE�V��wY�������ѯWZ ��6$`��h!�K���y�,�*�#�F�q�Cf}��4����b����V�E���x�X��nH,!�#�{u���{:�`���������4G�*���ī�w(��*��=�Я/� 2,�Q�͞<ee���}��sX�|��/S�3˵{�#{S����N=k������� "X��@���M��UNB�f���&��F8r�"�a���N�x�1P�aR�٬�qY:PX�X�(�]��vZ4%�Рz�����1��#�Ư-�C�]a���L�1xa�Q�W6`n"9	�� {�r�p�l$7����C�'�n0�TH��JG|�c2Oj���2š���FG_#�����\�K���^����|�҄�7@��}��=V�|>���fnm�2S� ]uY S���=�9E�+W��mr,��M��r_)^$V�
:�ˁZ���+Aݓ��G���w'l�5�N��NG�Q$���(N�[g��Nҍ�����+H�+լ���t�rzh�7�7]�+�Hٚp�p�*;��9�Ɖ������Y�qG}N��`�heq�������vŭH��@�(!�[���N��U����Tf~1n��#��
���v*�~���kb?�n�#aC�MPh�i��ō��k%o�Σ�/ꂄ�FW(C��@��}�I+C��~�#ubAn����}**!>T�[=I��r�+��EI1��i�c��C��5�"G����D0�`݀	�'NN�.Ͽ�FbOQ�8��$9qpb���:z^�	Y,1=TJ�s�o�����pb�� u��?�v�5�����ٞ�B�����$���X;A8�A#"|n�j/�ʯ�Q�+�u	��T��Z照E�(��^�\P\>j��F�%� �0Jى8[8���D�����m��Byh���,�4x��E������Vm��>�H�3&ռ_78\�
��]����� ��&N�i�ۖ"*��>D^a n[�<��4P����:g\�0l'��)��]�f�� �l�c7�&�X���<F�<>����DRʂ5���VhiՅ�CuZ�O:��~$&:)N�nr�:Wյ�j����M2/���'Q̙em�0O$�'z"Y !\��4 Ǭ��'\A��㑱-��`G5�RS�2����[��,׃�L�W���U*��ۓK2� �]�Y��f�Θ���u��@���kʱB��WE�&��p̐hn2!DW�K-�WZ�H�k�u ��f�����w��6��O57�F/�e��"R �+��΀�j�]�&n�H@ Thf6NP�O�X��w�w�sJ��KYe����T'�"zNA"�k,-�6v`eƉ�ȁI�pQYb@"$�Ql�<�������]XXǒ>�v�V�����	�=M��#:��j	�i��i/�r$��5��Z�{��'�к��.�u�, �����x�ca6!�0:b��Q�,�.9�Ƽ��*{��n�5r��CF4K+W!�e��:�(Vo~[���X��x�~X&�*� =�VI���p�����AQ!�uL~?Vy��ƞvX�<�no�¨D����w�ΗPN\�ه -��HE?H}�s@�]|�0���3�A��H	�qߛP���(3�qi	�b�M��M��>�;�I�:����R\*�]�����2��|��l�~e��-#֩��Tu4e���8�J�xN��mGִq1��|q@�V�>�_�-)��˞D��8���P��4��,T��Oy�i���B���N��B����/
M�z8+Hy���#я_�Δz�}m4�����F3�]�Ʋ��E�VQ8�άn�\s��s���JF{��芬529G�E�`?{�Sa��`F�D!�Ѫ�����/ i&�,�ZU�v�<��f����S=9e��K6���_���4���I���	D(�
�&�Cu�IP�X����E���OSz��@� �\�
��-�ʔ�9A8�guT�)R`�R:*�^b$7�%fD�άԼ�?�.�0�(C�hA�Ϳ`���4I����ZŨN#"Ii�e�S���\�hq���<��7K�0*��-W�|�؀�k�����j3rIڐj/cG:xO�,��`,O�\��6��YU#�¯'=x�u�G�����q(�jhSBI�hJ�2(�:�+�r�$�@���8y��r��c����^��!kR���J�	S,��d�m���]�X�mD�b���#JL<E�B2�6ȴ�+8���/�$�DMd�I�񒬼d8Dph i�~�:�1���	�H��{�Y7*V��uI?�"u�B"��4h{n�����"� ���M����Ȅ@Fki��,��L�\�N,.�2�R��K��u��S��:[i�O�a���h�x�qH�Y� k{"��C\��&�-�^؇<���_p2�-*z(�}��':aJk$Y�}ή�A9�/Ԋ=%� ��c{ W �IJ �I��-���x�8C	�h����b����0���)z!?3�LO�����Fç��ˉ$N_�M=%���TTCu�$��B8
g�N8IWi�p��X����jy�@V��'� �8�L�ʁ��Iq�i���%��q�"B�E�씹]�T#��זXf�<���;cq2�VRLp3U!�EYCj)�U���K���a�X��[�#�)�\��E3��I )8����{��^Pf�1c]=}�ݹ(8g$�U�=� �������{�̮�+<��6T9���;*wmf�����?"6,aa�dk~����e�&C
>�0��Z���o�M�y�%�H�d���V�0A-�̹#C5I8���? m���23w����[go�=u�pc���~N���y�C)���M�������6~@�&��*�_��Љ�����̿bn�hK�M   p�P��_1�s&�*tAK��;�%xJo\Ir�s��n}6<ҧ�j������H�ԲK�(��k�����R�
X*�!�^˭)��@���ɸV���A�<	Q��c��j�B��G�={4,3��<��o�TΒ���~]���ַ��������� �89^XG(���:vNbb!ºr��Z���Pn}����w��xUz	j`D�T� �XQ"��T:�Y}�_�=D���&��޻��񳼪r�4so����zweuY��'�b醙j,dn�b�l��F��|��zZ	ъ��X��94����ɘj&����C�elRZ��ct�b��}�G���[O,_�!���,����p8+�峱1F�PJ�fJ��1�������Oe ֞9�� �|`//�Ѵ�9�Z�ʶ�hGU>��m+l�h	^����9�,=�aU��3��)�6d'4{��`$�ݎ���8wX��;{o�Y^,�����?�R){�He���WB��) ˵B�{����~M�Djk����ԗ"g;jL�V�z�֑�i#���'�[������u� 0-Aɑ+Hb��� ����ѳD�WWߩ~�J��S��gNMʼ*�xh���V�$��eH�[�`����%_X<�Q���1��ǝ��e�S��
���� ã����)�)�f�/�ή<���J���UHz���LBj�$8����xT��v�өf�^W���4�%��G�f����T\�2Ѓ����۹��$�/`�w'YN1ezE��{��QJ{����𓛔��-2d��bG�!%��V��'��c���-R��.�IۧwC��J[���?�� K�8"���(�T<�}!�)ؓL�=�_������I/�� ����2pt����*1PJN	G���Z�q�ߩ�kv�m�o����v�J+5kj[�AQ*	�X�Ҁ1�b�?6E��L��)ƌ`6c��D)<@�+(F����^U����"�7mZ���M�� n=}I['�
�d���B�N��>1����z�%W˱������V��Mc}�����67r�D^j?>:����9@�v-��bf���mj��՛��g�k�����@�$���ڑ��h���^i���X�<�r*i�5��"��M�w���+���*+�Ý���)@ێ�?����ea$3]zC�}���h	������0������k��ջ��� �D}�@]
Ji�
�G�y�m��8VZZ�
v�",�r�"d�u�Bu3 ]N��B@���U��p��� s*����l�>��WQgU^}ĖB�:�v�)���.��yW0�n7�)��E�� � 5@ʿ��4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk���� C@��q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L�� /@п��U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM��"�砆�p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK   ƮCY�u�Q�"  &  /   images/9f4fed23-cdd1-4fb4-bbb7-c54436c6c6de.png�zwXS۶/ҋ��RC�H�@���DJ� !�^BQ�I�*E��H�� E @�)
��}������{�{����oe�5�o�9�o�9֘I��(ə����(u�5Lp�-��HJ��d��r�]ȼ��|��(��kxY97���v�K?K���H���L��»:UP^PG�� s�{(��t p'%�������:���36�8#AN@e�"J� 	�PHw_y�����+�(���T�j X��=}` YqaG111�,H�A�Y�H�I���K��KK��KHˋK�<���|���M4��9�I	����%/*(()���"*�D�$D%$�qa� ?(J�×�/0_G����p�u���S�T�w�O��2��L��ET\DL�/(�o�W-�ű�_#QP�:9�����q��%'GQ�;	����a���z�z�y��z�7��n�wK���g[�ȿѾ~�~�3��5��z��8�4pfrWdɫ{"�|`��8����
�����Q���C�A���H�	1���)������W23���+���(�����?�����&�j�����K^���i�N^+b���	IyiYyi��br�bb���{:����K����ؿ@q�8A���G�������s����D�<\���'G���n`���먫�x:��qZ0�C����+���u<|���0% N"�;�KJ�88�ʈ��de���` a&#,�9�9��KJ���_����*�������7�4u�_�J.h҆��y���tMa�޹���<��Q��9��������+�����|=���>05���8��& !)"�ׇ:�=�$ust�z��p�U(�sG�?=�w�E�-a�%�e�?�%`���)�S�KЃk����8>�h�AP9����>��u���e�@��Rf�v���qe�N��iƎ�7y[$W�>�p������It��F���MX��\!ȧ��7B=��#%p,�c�Fs����'
1���~f���NZ&��H�s�� �	u0O���R��`���	L�پ3�Y��z���o@��tr&31�m�Ĺ�oAX�V�0(TμtL?6)����oM0)����F����G�1�M�g�0ؚ�گ/��,2���؎*���<tQ�܈�vC3�]_ָ��Wn<ٙVJ�ҥ������a||�}_]��SV�Y
�	ܥ���ʿ- @�{"r�~3�N��,��m��m%ry,�|:��V��))G��w|���e#,��xM�ᯠ�בu�T�8K��-!'ߢ>g�
��A	ԡg��b�0��l�.ވ�"���:�8�m('���x{����qQ�~��j;��2�!no��CU�O�	<m�~�)\�U���ƾ�w��C�� �F���B.��ڽ5.��߼{]p|��W���m�`�H�������;jfv��4�[�������T�$g(��OX^�4QG'��LK�bP�
�g�Q�s�
����B�][�~{LEv��W���t�y�V,�)�8��1M]��PM7�y������+#�ݴƙn��=�&['1��-r����C�G��ޫq��ö������c�g�aq8�k�}��
���F%�`{ycF�8D�ԧ	FR�����-�3]ي9�ׇ���W��j2�컑�ґ�����u���&&F�-:M��N����wB"'�w}Osp*(���$K����?F���<�c&NӢj���n%@��w�b��ڎ�Rj`y�L����Z<�L4��,���֐��Ţmy�V?
N܀�&Q�����Xqj��+�:�r+��`A0.@��1�w�"��)���X��7	�v<f���S�h��i�V��J=}�����d�uin8}�掳��췹+ݨ�!^�N��4�����Y��&E}I��˸Rr��wӣt��1�����72�����ҡ,����_)H�$V܌Npɧ�'�tw�a}C�:>`_��j�?0���(�#�bzr!�X��F�P��bD�|�ݣ��MT�r�Oњ������ߴ�k�o"]!��A�tE�ʱ���~��i�8|g5ܑ�D$ �trZ'؂=����3��O�����2��-vn�r���^׿ҳ����	������B�R�!y��o)P=TQ�c����*M��N�<k��EMDT���}��~S�( �Kms��j�2����8��F,�G,V���j�Хld���H1�+d���`8o��������:�)K
�a^[�XT۶uO��D��1�v����*��7��Fg�{��k��"Z�4��
p{�D^6�t>;U���3������r�%r�UU)s���J[YY]���
�&�\��T?gY� p>������64ܶxs��p̰�)��V�L#�=gzbb"*g.@k*�uq!�]��B� �k��ZKwD.V��A�ì�CzY�sVi�l�8ã��4<L�w?,E�Z|�����z��4��.1G$Ǒ{Ě�M��b����B�I��4��?n�5�+���(v����al��I�^�����4�Hr\~��.9���3�#]���/.r���^i����5d�/r{Tbd�� C�n����KǍ�U��9kC�z��Ç�^}
�l'���I�[��q�ڂ��^0?1I����hͿ�,��	�m�6-�����w��W{�R���1C�dtO틥��UUO>���.�|�'XP��5�}�&?AA�FB11����%+[�tla�������S?MZs�}���R����-�i��$S����4ת��P (����-�c�A}�\�Y��ݷ;�CZZZ��\I�!�詼#��%����=;吝�%��Y��S�l�SVèF��e�>������u��ZJ�$g�;��Ԍ�<��X�ԷDv�yWd����(&�9���i����}8�!|�̦p��Y���r�A(��:��d0� ����"��Rq+u\W*��=NE6A����|��X�sm����r���M%3�yx5�h�u���������vYn����T<���|�(�kb�7P?�`}�C�ϳ���®��_|��ќ��Ei���R.C��CY+tܐ����V�+Vֶ���/<�9��T��񽙏�E��˳XlD� ^S�F�~6ӽ&�d֛����z��u�>C��a;�ikR��� ^q�CNF0�L���V���/��-PF [ ����9N�G��M_)� ׾h���A����[*���u��f�I����s��{��^�J�vU��U���Ѫ3g�`y�b�#`f��a����P�Q������.���HH,ԅX෼�|�u�\�Is+��؞�E����4��\��]A��r9z:7 OW�Tz��Vx��Y5�ύ�f�.����P�b���1���P��M��qZ[�\����5�gkEZ���[�A4L�������h$���$�IA"��;��B7�Z���<��������ý`�F8[�����֡*��>��l"n*�T4�3��\�(V��L��ԇG�~�/9���T��{�a,e��,��<7r�s�ҟ��5PGj`$g��3\=#y�6B����C�(����x��Ҭ���X���*P.����#n( ��M\�zL������L���qcZ,3����7B����f�ucXd��)���
��S@�}�*1/���'�<"�W��08]��B�4>~i0I��*�h�Z�ҧ�+wcΖb$��j7I��.���p&ବ]�`��w��и{�@G9�[����Ac
ڌ�BdҐ��17����mk�+�I|�iB��	��ڰ��K�[�)覘x
��]U���^0r�ׂ"j�)A�����E��^�|b����e�8�wf���UL<��VR��Z*�[mCS�������{%��9�Hqڇ�D�es�l�e�WD�[ʘ�6i%��.�"�B[h}i+�u�P~��/��(:d��������ϞZ�7�}[c��>f�΍��6�!"z��y��+��u��9���V�p��;�����y����\	����מ!`����B;����_���Qi�t#y$���I�rަ�4%�kt���:���')6���h�a��*ǽ�>i�������j��:od��*�q�D���
@XM>&v��0�!�)��%��׾�wAޮ�̎���**����hkB�Ѧ)�x��/9e..�,D����~"3;<�d�O������F?W�8�����'T�(t0L3��[~Ov2*JMIӸ�̈́�>cy��bj�Iy**�`�Us[Y�|��ME��Ô_��B�<
���c��7XB�㊨x��$n��Z�㖧Hv��",ܻ��˿��0�#f����l�k��(L�Y�W�ѫ��cޮ���\�q����T��VONŭ�6�T*������w�֭}Y���:98
=�!~h�I �� }9v�)�����̩��c3Fހ���߳�'��h��b���9�y���Y�V	+0eO�!�y�»����l�<氌����f��>VJB�-��A�V`�h.s�r�f�|{�u��r4[�+�#�şͣ���zVI8�6?��� �U�[����uj������G,R�'�vp0ܷ"s<_����W�͜��B�;#�a�aw��k2Ebg�ƻ/$�����{]�<|��c����|a�N`"�\�]��O�\�2#�o��/²���$�����x�30�#lB\kw�W�O�LG�~�I?��g>��k���7����jM�ȩ���Q_�.d�r�x��������5=�vY�%�����]�Qשd3N]0c���` �s��C2����/U� F�)��]Tf�~��b4���ȱ����pȒ���_�;c4��xB��sB�oL�Z��*o�C��I�.3g��2�e���"�{�9/�� V��&:�M$3�[���"�G�+����Q�n^��Lk��uܞ�:~���h˯��J�d�יɉ���[g��ׇ8�mT�%�I�hE������|�N�J8�#�Scc/��'��M�Q�=���n����އ�oo�r��#��ϲBO?D���+/�\J�]k�U�7ڔ|ů^H�v��.�W*�H�NY��T�t�һqN�VO+�Gi.nk�Է��V����si�44,]�[߀[oI�y�i���qF��
�%��y.��>��I��̃�2�d��Qt�+tX�7d�7��5=\2��q�;�[�[����m�ǒ�˵�PIV:��YWz����C6�\�f�������U�E\�苋���-�l�Nl�T^�'��ƗD�����#�H���J���,I{���7 ���g����]�rŗE�7���O�;��JKK+8��<ѡq��Z������^6�!m:QKT|�m����s������I5��6Sa)a �R����� �xI��q��8
y� j1���F�.U*�f���\�1��%Fޤ+kk���I!�O��7Q.�����D�Q\�����z��J�2���]9t�3�,mHN�:r�ź!t��'�� 	l��)�RN?Q�׍�s����WS������y�OϾ?�T��)N�S1�M��>;�
�dW�y���C��^���ާ��ΐРWj$�5,�'�2��[(/u��)02� �Il'-�!�j� �7�w!۝�h�۷;���O/Q4���v�"��]U�ƍ��j:N´��6dӶ]�F�F�51t�\�jM�4�����G�3�6(���pB���lf�����U>whӽ\�B����+ܗX��j�3cg� ������֍�)%�K�D�3�Do,��ҋ�x�	��d�I�x���b��|�+�����V~������Ri�j}���Y#B+�,s�9JPH=]㝊����2Y����_'/�Z�HBIH;a�Fj1�Y��T9���'�{����#w��E%޴g<d�� ��w56ʾ�����2�&�<?�ɜ��64���?��~��z<0���}DMfތ?s,L��$�#���;�5Ǿ�W�&6��#M�%Ƙ	Z'�Įn��z����F��BL�����|��$ �\�t��Y9�! \r��� �Wٶޔ����R���!���`��5ns��"��:/���3�O�CE��5q��T�Ѝ�
���T�3��*~��K8Y���	]>��7���X\�l���=غ�3�6`���X8��$.nI��ۤ+7Ӵ��j��Ȳ2��#fD�z��&�����:��ɗM�tK����<��}'/�zq�Q'��_>��_�W��}ͤ�����AP�F���=<����]Fȉ�����T#�#K>�ҥ�W�^���}`�(�1�HK��u��_�*&��O��x5���N3�8l��h�a��FK5���֓��;g��I���MY���B-�䨐�����&�@<x/v
zǑ��C�Pu�z�:�϶�'[#E�n�D?t�W�n���é�"E	�c�0�ց۫t&�k�o3�)L��8�]��z��#|��ߌ��\�3�`C���v���%��E���G�/��ށF�g?'*l_/���z=�"�L���[�S��_�]M�O5xj���W�4'L�\
�|'YՐ2ۂ���Rl'^���{p�6�8z�At2jb��h�|N��+((�2�ۺvQS�デ=�Ͼ7��tŔ�yW��q��%�sk[�Bf-�>Q�=&qif�u�=�����U��:A���]d���m(�RD{��z��g6�9��R]QyWϬQ�U)��p��pÂj3)�d�W�8�}r��N��Ni���(��oM����� K}�M��Y���a$����P}���0q*��� ��|��A���R��=�d�'�������Eo��F�fSe����̹	-�����ɍ̲l�n�RT<2���E��2io�x�6/��?q�f{*}�bU>bD� ������� �G��K�)��6�S�֩�����Ln��z��
M��s��^�&d)]}�L 9�u��S�T
?���ӳ�|.ݳh��$�tr����Ȥ�?�گ��E�=��˝���S|����Ɇ82X%�TƳhlG����	�;�}$N${�ӧP^P��&� 9��c-贠����3Ao����e�g���PEƼP�I�i`Da�����:���a_q1H������xS0���E
	w]�~�O�8��Vu��h�?�i�)���H����_��ԭ�C�+}��H�Ѿ�DXd�`�>��&*�_a��ި[_�؛��iO-ڤ4no�o9����u��f���-�Ǣ[.2O�"3�iA2�򛙯�γ:�)P�4���G�YB�#�8<���?�	��.�n�E�%�i��Xۮ��ҷZ&���v?b�~uI����90���eb�ԛ�ٖ�Ơ�)���t�{�̽�64��w�O�[Af7� ����>&p�8���ڿ<]� ���X���;Y�E�U�'�}F�>��2c�>m+�a��닅�ݡ����1�h�n�w�U�"6~�@�00"d��Df/��p!���V�z�b��x�}C��Bzg���\8�G��ϰ��%�){]*�p�@�4X*��C�˾�t&�?W-�E��Λ�N�OXh9�~8�;{h~�����Y4/��Aa���w��B���9��o{E�H�XЦ��m~��=؆�PjuI�.���u��{RSn����~j}�iAh��u��?c�ēõ������E},���h�Kjfn�g�mKDqO���I��kA�K(wNL�Z	-�R�^��
6���G/a��HG�������ٍ�/E/�^��[3��N�Xb �ڼ�g�tqR�y+���>���X���E�#���1����ӞD�J,x�s�����(S�U�{Hp�����:����M]�E2�����e�[
s׉�F�آ�/����wb��nNW*��u�$Hh�S;O2���dp�����ರ�뤃�����~+�w�����r��FRI�a�8�)��Pr�����[�}k'�3������U�?NX2�Xï�v��'��H{V�VV�Vz>��J�]鶵S��T�zWQ/�&u��I��&]4�xe�rT�53�.�Mh0�� �o*�}�|���d̬0��]h�p`���վ�ܻR!DRU����!b�F�������I[|��D���e�����h��Tч�`q�*�^hP�1T�|�S��H<ق��$u��Zj�l�+����f�ɶX>�Ņ&�~۞청��ZM������ڠ}[���Y%v��_��o/lx�8v;�{Q��cKQi]fA��Y;�IE�ֲL�������j���!�����U���55Ɇ&r4�?�u����L�ro�!H�V����~�G�ʴ����ajjM���C���Y���ީ�K���ׄaaa�$6�k�x�q���R��S_��L=�w��������ӵS�|.��W�ɉI�"[�@l�'|=�VԦ�q��Y�?X�(����Ti���ÃDM�Ɨ�?h��q톸��������C�T:���*�K��Ξ)�?����ښ�|�"�>��el�}rt��Gn�� tQ�eU&e?ol=�2�{sdn���8?���8�^����/QA��W��L{?n���D...?��to����}�/kF�UWW�l��
D�)�%iUn��o�/\.�˭�f)���%!���)� ���۞%������vHa�E_a���3��Y]�|��KM5+��p�r4SZ�Ǝz��r�	�6��Ӱ���,��){5g�r�	��0��w�ј��?�.�M�ύ�Y�1��NҎ�Y�~S�9Ufj���]�gKG�@��>�? PK   �v�X��C�N  I  /   images/bbeacf7b-7208-4b04-b839-dc1aa989c418.pngI��PNG

   IHDR   d   S   i��A   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  �IDATx���U�u��0<��y#�W|E�b�M�5V��6�������Sc�hMl�1I�G���51jbk5IU���F06A"UE�	�0�83�c�a�������s�=�{��~]߷�{�9���^{=����7`��ɦ��ǿT+8Qp���
{w򅱬��1���z�B��O?$8=����8��}����8<�}�1A��'�s�ۥ��r����C���O��ÇM�~��._�
��54���u~www�D�
t����wK 8�Np�`�`���"�>����0�mۛ�~�3v�	�_���r�u��R��3\�g&�@]]������_9��Ѓf!=j|I�E�u��	6K��%��� 8Dp��$�Y��
��#86���F�7hР�8y'΁�	絋��'�U������uMxQ�Cͤ���ꊈ4��^&���1v���C[��@�[p��s�fm �s��y���f������Q;!�rK`\ ���͡C���&�ǂ�'k�ȭi���y���}������g"
� b����|Bp�I�?f�l-8��C�S���b��竂���/c�}�������L�7��O�3����\�`~����N�jC��+��rD��$��f�w�Q�gq��H�~k7v�R���XL�so0V� �]�q��e�o��]"ߗ
�zX	��~0�&}� �q��'�5�S�52+AJ
�`���r`~'E	hY�d��'�%����K��p!�"���D�(��?%�Y�q>#���%�	����-HDc��S�uttDc�Qv���� ���@2�<��Cs0$
���*��4n�\�P����N�/����
n�5c�!S� !�pH}���6?%���|�Up�_X��0�>1�eT�;�H��~�=dȐh��L@�3�>�`���zfWða�v�{�ƍ�˭Ok�1��36g� T;�T�4�*�E�{�7+��J���I?�I�����	��P�R��*���ݣG��b^-?뛛�omii�$�8/�3�˂�͏$.��#��0�,�	�A�@����1��O��q 1mY�bOVE<��t�҆�����,!�b�U���ۯ*c��D�@�Ϗ)S��-[��k��Mu���Qx��#��F��!��\Ey�T%��BL��|�c`�|�-�lr��?'��`S�=q�����8S���/�D�rW
�,�wq�)�,P�X��3���X/�{3�A��1.4�X}B�,Vtm۶M�Yp��%t�.�r"R-(��_�Q~�+x\X^��<P��`��:{`mt�n�{���}F� -��3�}�TF�Ǔn̛7���է�P7jԨ�{������v�?q0|�y�*�!��|�`��=\�x�9�����C)f0��0I��X ?�/,X������4�]xekk��q^����	FO�
A�4�� �#� �ϭ��"�������3g�M�6�nz�f��Y�S����2nܸ!��A�뽂��b�e�p���-�8DT���4�'YEWE�E�#0��&oV����� ��9�FP��E�������f":��y��k@Q��B,B|��	��o֊�F9��]$U�*���lM����O�� ��ޒRn{���Ks>|�� %Q���o�䎎�C2����P����a�cC�K�^�UAQE,�G�����8P-��a��w��%�MNb<.3|�����4����|�'�\&�xF��V�>*�*�����ͥ�^�+
��x������5/��r���2p�0�	�qG�2{�V*��	&���/��M4�ս�bM	w|9�
��]�W��`�/�ҠAtQ�a�k{<�%�@TUCo��"��]�n�{�tV�E,(O�M����E�"!J�z�!,(�����2T���@���I�,�K
����MG�	��̾��ZU�����<y���s�obz�9��2]@��Sf��?��}�m߾�O�/���Z"��j���Cc�"�M��IVWn�0�@l0VnF�=��E���Y�_"��&a�4'\&��W���{�d o�s�|��Y��_��kiiQ�L?N��FV �&V3�׋IAH�J����������H/"�;Y�F13��<���2�mӦMC���"�f�PF����i��7���755�?Q��h'�z�޿���5�d��l�^}����I�&�k�@8B^�7�����X�a!s��':�h���뎝;w*q�ٻf�?� z�5� [��o7v�J�J���_�=����4��x�c�E�Z*�#�r����666�'��Ῐ�7����`�}2�|3�:�g��S� �6���g)a12+a�?2v-39O蜥^�~UpP����o׆�5 �I�f���} �����}���YwY@	��TWI}ɵ32V5��D�"��s�<?!$@�Θ`�L:�b�]�
!��P��X�gJH�~)&�_�㵒L�
�hӀ4 ,�>�4�n^������[u�@�_�%��,j��9�L�:��͛7�Q6����e��@���u���* i�������U��"!� �K�ڵ�T 
��M�6��-�2��.�p	6:��mG�9GO0vB�O*�� *C��]xX�p�8l���w�c�-�e���r�D��1�|f��*��f�	
W]ƿ���������zIN�GB�y��+���lv�X��&�yR������$3�*��s?ق�Gj���M��a,�l;׸��N��!T6�X+���ٕ�^�QD
��B.�����^��!$����;�i!��g���A������L�X�%+����E�(�=�P�̒�r�X�&�B�u�$�����Դ_���ls샆�p�Dd|b�D1��������OV���9��e���ث�Ʀp��
ΪnY`�M`b�56-	O���'��� A����J�"	�Q-B��!q)DY#ˍe���fo�����I��!��W8C��VWlJT�t��y������-��
��Xfv'$B�c������u�<"qr�=���[$�r�b2�rc��z���"�M���2y�VT�9��6lX���w�G��39 JL3f�Y�zu���YZ]Ie�z��s��5���2�{SA;����BC�i����on�ԩSu	7�ayCB���Ŧ �HWID�rVqf}�A�ys�M^����S���	10]��1�F���PF��ɚ	Y���M-G�V$�j��B�e�Tͼ�{V%�� B�g8d;��4����J"�qH8(Z�цH�5G�� W������<�C��è�<;$�#H��ˍ=���IKͱ�]�:��fAG�śBd������@D���At��'v�9��~���o���Y��_0v� �.�"��W�c��Gc��Z�`�w��!��,��+�� ';˅,B8�M1�).)����f_ɇ����g�!i���K��'	 �r�o�W���dEh�D� Ib�ƾ�c	�{*�8��������z\�����i7��3?cB�`��=����I@�P̕����$e�j�%��"Z�LG�,.S���+zJ�b�F�Sɣ�Fp@1�m.F��9J�am1��r��$9`a@�����⸩���z^��֮]۫`@�\���lm^@��s���M�ِE�[ӀX�g�+T� g��������c�ql�z�?��=�q�6`�)�ω�`��z�^�\�5�ё��Ϧ�%����EB62�l�o�z�8����n�EI������VnWR/���*�������ȭwĈ��N��UQ�ó����*�JJ��Y͌�L����E9bx��:2��,"�p�}��� ±y�L��o��� �X��E��PS9�TM��ⴂE	5ֻٰ�.�R�ܪ�r�#����p.����~z����:t�۷o%��XeX1i&9��F�'nӏ;��	�ۄ�?[I��ِlV:.�`Q���XXQ��q�)�DIN<�%-71<?dȐ�tvv;R����V��B!���0駶8�a��O����y\�	v
<��p%�C{4_�L�Ę;wn�\FQ#F�@��r[Ȇ|�7�#577�ٳgG�ۺu���A�e�g�X������\�2~�x�6�Z)�9�\c�_�(��L��L�� ����u�dV���;�q�t�4���K����E��q�~�)�&�Q���!�3�Mr�����w�!)w�1��fp��?	@R::r����>��� b���e����(Z�9g�+���,�P�F��q��utJ��8�m���vD�s!�ľ�^*�C�Y�'Z�.ܒ9�FS�@�Q	!7A�%Rcu�礡rއ� f>J�"��H��y XE*ǲ����y�G�<�_�7�\c<x��H��F�]?hР�ك��I�
�V��0�Yed�K�"��t�*�@t�e��G��'��=R��]r�V���+����l�C�� v��p�"�\l��U������Q�w7:nY���K(�3^X��&8�w��{R��)XR�]"�Q>Sk���o ��Y�����d=�"~�w�H���/w655�����Fyk�u���!�*�`�$(���<sD��$Q�,i"xL��+��2T���J	�?K/-�1��	��lժU*�XGG�ÊA�����-_4V���`�RVO�. �"�a�g<)��G���{!
l}���M/R�3�B@�UI��u���� K�;` ����9;�0�~L��K� �〔����}��n����5����!r�r������Y͌#
�������ߩ����J��(�/1BQU�KJI*rgk��yԨ�!]]}䎞���<Y��5v��PI��`;3��2���pPduA���2����E8�pv�=GV�e��ұ�*͓�r#J�����ڶ��/��/j��o +F'N�Â��ޒ���t�ia�� 9�!�� )����刣=@y�Z��=��v3�>�_*3�N�eVF�hA5|�BHƜ1N�a�EoE8��g�k83Ɣ�7���[]��_�>X���o{^`v�t���]I�>�Cp`��Nu�ݙ��4���	�Ń߰{�nD��~%pF�7�a̱�鐾Lk����+����~B�|Ѓ�P�QP����]�CX3��y�$��ve���YQ�:�Y&P�~A��1>���K�3@��Uro�|_V�����!�Dx��%����d����55�B�ڤwM%3��B��*��]��v:��ń���th��)� 'e9�&��{D�%��,�*�G� 7�����zC�I_�]*�Dw�9|��Ƭ�x���Ms��Ɖ��W/����4
1Ȓ��݄(�<ĩB��;d9����b���d�x�4�����m۶�<s�̗:::NOz=�B���LT"�h2�<�?��pa���p���`89�>wn�K�"�-q�!�sF������b�8��C�Nj;v�g�3N�ed���a�{GD�bq�a�{��:��}R���#}J<�(y:����Mc�B���:b��$	;�#C�Pw����j��A�gI�G��&�,�mH�ަ�B
E7���I�
�����I(%X��g$��i��i@p�/�!�p�W�=���1���u�&�����m�__`9A��)�:�����jڪ���C�ꦯ~J{�E&O]de����=�S���eM�3{�}M����Ʀ���nu�(#�&����� ! i?��ܻ�y$���#t���ߥ��qqi'(�e���{�[�|��;�3G_&pyJ�ǩk�����U�Y����u ����+4
]�Hð��`q
{F9�]��}�ɞ�"�(L\�
����?g%�9�¯�K�T�Ǝ��w�� l}�t�H)���l��kG�v,i"��G؃��w8��>���$LF�~��#Jc7���r�.A�ϥ/݌���PPV���KAB=�_�%�+T����Z�n�,�rѓ���1�6�Db��2��GXRE$�e��Z��:�5��:Y�_�K�����}�Gd�b�"�������,�P٪��M Xn�C�9~A�<J���z^:���ۢ	��~�_ �p�,4eN��3�}��}ǔer��C�<A��GD��x!z�Nk��HE`��3o�8�4�M ���A��_��k�=d�8"%sB�[pT��?O�@g ��o�3���.8�b�W    IEND�B`�PK   �yDYZ���  {X     jsons/user_defined.json�\mo�8�+�?�����~Kc�!@�N.8`,(�j8�W�SE�����v#����݁͗J����g4#��6Z~��ѻ�j��ߜ/�ڻ���ٷ���� �pF`�b�wC�w�~{ݸ�Oݹ��[FaHa��S�~�!������|T9���\0d�����!c�@�J)�6'��i��M���ë�|��+޻e��[��~Q��|��w��mU�6��3�Dr61W�2��u\�\%�,�ן༪h��I��
�#�w�
/�1�U^kx����'��h�o��࿳�
[|�pt^�Wuٌ�}ի�q������f��@`�&��M�/�c&#Z���}UW���W�W�n�V`�N7�YT����"3 %��1�w7�Z\��禅�_�7���N`l���0<	�sB×v������x��p����A|���(|:��
�8x>/�:~��a�e �DF�>������_]�7*�>zЀ	 �G0��
�P� J�-�$L�!�,��B"�Dg�>d!$c""-��0SIH�DF[dҾ���&���}1˓C�p;���<�"?��Y�L�1N��/f���X�و��,��E��a�Ҿ����s����5 �O���x��c5&���*������W��+{��(hX���� �C�b?����9���ZH�Ѹj��
r�㺪��t>_�Z�ﰫm�]V��s��6�j��^4�YL�c�(��)���Pd�Hy.��z�W�:�1���^�
��b
iONZ��p��u4U�iL-�G����s�t))��	�t�#3�T[�I!=�աP�*udJ�u�t:�jyB���1�7��T�q��7��E���������������������������������������������ܻ��À�������ռ����74�Y-���7�{qcMj�#�$H)c.G���S�	\Q�b'Zil-r�Y=��� ��`�0/��c�Q�,��]���j^�H��93��Xu���Eu�C�0���;��nh֙2��nԐox�>H�~(C2c�zA?v�"��Ϊ:���&�p�HЏݨH?.�*�Ϟ�$���RU��Ѿ���g��|O_�^�@.6��6*{�װ�lg�n���.C8�/���|��/!�o=�d�P-�������Z�zͶ.�C�l�*m�\���3{�lٮ���U�V�9��ϻ��N(�x���Ý�$Y�r���=�ҙ�E��n��H�])w�ܕrW�])w�ܕrW�]W��F�3ظ��a�Ҷ����ӘfX)�<��K��9C9��)��4F</�d2�R�;����"[f�T�䴟�<��ݿC���C'>��&�����g������MlH�2�q��m~����4�� O(���Dڟû��|�X(?<��?�w� �bs~:��ܟ��fk�r�)A���0�ϔ�O�� `�q��} �?�w�@f�G��W��Ԉx��۟���������-��������K�K��iv��%�,�ُ��h �/�~lz������Ï�n!XG�30���2���}Գ�����
���L� �fz6�^=����tz5��%�m3kf���ja�T���,�1��"�`�$���T���%U-�jIUK�ZRՒ��T���%U-�jIUK�ZRՒ��T��7V-��jy��R-�ϣ��ب�h�����(/E��қ���v�O�����#M�E\	�,7��Bʲ�F)Z���SzE��TU��"�0�&��P�e��c�I�Ύ������)�TO�������\S��;�P�A��9��\�Bp�d�'�&�&�&�&��/2����{���*k�J�S�#�A@d�-���b��<���>���tkc�ÈӲ@��/���ཱུ1y�mQ�)�5�9�if�+��F����kc(�$��YP���*���O�_�L��9e,Ji���?�����/ia�q���!�������PK
   �yDY�#UםN  2�                  cirkitFile.jsonPK
   [x�X ���s� �� /             �N  images/14933c3b-4ba2-45e6-999d-97e61a94bbca.pngPK
   �yDY��� 1� /             � images/1e4fa634-4e77-4d97-9022-ac13a26749b2.pngPK
   �yDY�TV�w'  r'  /             � images/3b67e01d-51b5-44ff-99f9-fc90dd618da0.pngPK
   [x�X��"�IY eY /             pD images/42bd9711-1b72-4047-a3d8-ad461b8cf403.pngPK
   �yDY\��䓝 Wt /             �	 images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.pngPK
   ƮCY5��<O  g  /             �; images/4c6ee15b-826a-4754-a49c-440dc66ff58a.pngPK
   �v�X�}��k �) /             �U images/5b84a191-11d0-42fc-8d11-d4f69521b0c4.pngPK
   �yDY���  �  /             :u images/5d57974f-fced-4f10-a93b-7d150e366d9f.pngPK
   �x�X��/F��  ��  /             q� images/8278d802-2c3e-4ab9-9a04-8028f624633c.pngPK
   �x�X�ة� � /             r� images/8d398a91-1a51-4737-8347-b2d4588b3940.pngPK
   ƮCY�u�Q�"  &  /             e� images/9f4fed23-cdd1-4fb4-bbb7-c54436c6c6de.pngPK
   �v�X��C�N  I  /             �� images/bbeacf7b-7208-4b04-b839-dc1aa989c418.pngPK
   �yDYZ���  {X               '� jsons/user_defined.jsonPK      �  �   